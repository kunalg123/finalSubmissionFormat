VBGP v/s VDD [2V - 4V ] @ RL=100 Mega ohms
M1 3 2 1 1 pfet W=wp L=ll
M2 2 2 1 1 pfet W=wp L=ll
M3 vref 2 1 1 pfet W=wp L=ll
M4 3 3 4 0 nfet W=wn L=ll
M5 2 3 5 0 nfet W=wn L=ll

D1 4 0 PNPDIODE
R1 5 6 9K
D2 6 0 PNPDIODE 8
R2 vref 7 82K
D3 7 0 PNPDIODE 8

M9 a 2 1 1 pfet W=10U L=5U
M10 3 a 2 1 pfet W=8U L=1U
M11 a a b 0 nfet W=1U L=3u
M12 b b c 0 nfet W=1U L=3u
M13 c c 0 0 nfet W=1U L=3U



Rl vref 0 100MEG
Cl vref 0 50pF
.param wp=12U wn=8U ll=5U

Vdd 1 0 3.3V

.dc temp -40 140 1
.include osu_018.lib
.model PNPDIODE D is=1e-18 n=1
.control
run
plot V(vref)
.endc
.end


