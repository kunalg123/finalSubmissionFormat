magic
tech scmos
timestamp 1594279047
<< nwell >>
rect -104 175 131 418
rect -15 -289 131 175
<< psubstratepcontact >>
rect -156 -767 -120 -721
rect -44 -767 -8 -721
rect 61 -767 97 -721
rect 165 -767 201 -721
rect 266 -767 302 -721
rect 382 -767 418 -721
<< nsubstratencontact >>
rect -97 371 -73 405
rect -23 371 1 405
rect 51 371 75 405
rect 104 371 128 405
rect 38 -487 58 -481
rect 38 -687 58 -681
<< polysilicon >>
rect -88 346 63 357
rect 73 346 115 357
rect -88 329 -78 346
rect 1 329 11 346
rect 53 329 63 346
rect 105 329 115 346
rect -45 187 -37 204
rect -69 179 -37 187
rect -46 15 64 25
rect 72 15 115 25
rect 1 -2 11 15
rect 53 -2 63 15
rect 105 -2 115 15
rect 1 -305 12 -295
rect 20 -305 63 -295
rect 1 -316 11 -305
rect 53 -316 63 -305
<< polycontact >>
rect 63 346 73 357
rect -77 179 -69 187
rect -53 15 -46 25
rect 64 15 72 25
rect 12 -305 20 -295
<< metal1 >>
rect -104 371 -97 405
rect -73 371 -23 405
rect 1 371 51 405
rect 75 371 104 405
rect 128 371 131 405
rect -97 326 -89 371
rect -8 329 0 371
rect 44 329 52 371
rect 64 327 72 346
rect 96 329 104 371
rect -77 187 -69 210
rect -77 172 -69 179
rect -171 -721 -157 111
rect -53 25 -46 208
rect -36 -295 -29 207
rect 12 36 20 43
rect 64 38 72 44
rect 116 38 124 43
rect -8 28 20 36
rect 44 29 72 38
rect 96 30 124 38
rect -8 0 0 28
rect 44 -2 52 29
rect 64 -2 72 15
rect 96 -2 104 30
rect 12 -295 20 -285
rect -36 -305 12 -295
rect 12 -316 20 -305
rect 64 -317 72 -283
rect -8 -486 0 -462
rect 44 -481 52 -462
rect 116 -487 124 -286
rect 352 -669 372 -650
rect 38 -691 58 -687
rect -171 -767 -156 -721
rect -120 -767 -44 -721
rect -8 -767 61 -721
rect 97 -767 165 -721
rect 201 -767 266 -721
rect 302 -767 382 -721
<< pseudo_rnwell >>
rect 37 -481 59 -480
rect 37 -687 38 -481
rect 58 -687 59 -481
rect 37 -688 59 -687
<< rnwell >>
rect 38 -681 58 -487
use n1  n1_1
timestamp 1594253749
transform 1 0 44 0 1 -459
box -1 -3 29 143
use n1  n1_0
timestamp 1594253749
transform 1 0 -8 0 1 -459
box -1 -3 29 143
use r  r_0
timestamp 1594278423
transform 1 0 72 0 1 0
box 37 -682 301 -480
use p1  p1_4
timestamp 1594254441
transform 1 0 53 0 1 -283
box -16 -6 26 286
use p1  p1_3
timestamp 1594254441
transform 1 0 1 0 1 -283
box -16 -6 26 286
use p1  p1_5
timestamp 1594254441
transform 1 0 105 0 1 -283
box -16 -6 26 286
use m_l  m_l_0
timestamp 1594246348
transform 1 0 323 0 1 136
box -497 -34 -387 36
use p1  p1_1
timestamp 1594254441
transform 1 0 53 0 1 46
box -16 -6 26 286
use p1  p1_0
timestamp 1594254441
transform 1 0 1 0 1 46
box -16 -6 26 286
use p1  p1_2
timestamp 1594254441
transform 1 0 105 0 1 46
box -16 -6 26 286
use su1  su1_0
timestamp 1594254037
transform 1 0 -89 0 1 207
box -15 -7 27 125
use su2  su2_0
timestamp 1594254199
transform 1 0 -53 0 1 206
box -6 -6 30 126
<< labels >>
rlabel polysilicon 6 341 6 341 1 2
rlabel polysilicon 56 19 56 19 1 4
rlabel nsubstratencontact -5 390 -5 390 1 1
rlabel metal1 -4 10 -4 10 1 3
rlabel space -74 135 -74 136 1 a
rlabel polysilicon -61 182 -61 184 1 a
rlabel metal1 102 33 102 33 1 5
rlabel polysilicon 31 -299 31 -299 1 6
rlabel metal1 47 -475 47 -475 1 8
rlabel metal1 -4 -477 -4 -477 1 7
rlabel metal1 48 -689 48 -689 1 9
rlabel metal1 120 -307 120 -307 1 vref
rlabel metal1 360 -665 360 -665 1 10
rlabel metal1 111 -754 111 -754 1 0
<< end >>
