magic
tech scmos
timestamp 1594123059
<< nwell >>
rect -526 218 -354 311
rect -526 78 -353 218
rect -263 98 -173 311
rect -83 58 87 311
rect 177 58 347 311
rect 437 58 607 311
<< ntransistor >>
rect -477 -17 -467 13
rect -447 -17 -437 13
rect -417 -17 -407 13
rect -23 -91 27 -11
rect 237 -91 287 -11
<< ptransistor >>
rect -463 98 -413 198
rect -223 118 -213 198
rect -23 78 27 198
rect 237 78 287 198
rect 497 78 547 198
<< ndiffusion >>
rect -497 5 -494 13
rect -480 5 -477 13
rect -497 -9 -477 5
rect -497 -17 -494 -9
rect -480 -17 -477 -9
rect -467 5 -464 13
rect -450 5 -447 13
rect -467 -9 -447 5
rect -467 -17 -464 -9
rect -450 -17 -447 -9
rect -437 5 -434 13
rect -420 5 -417 13
rect -437 -9 -417 5
rect -437 -17 -434 -9
rect -420 -17 -417 -9
rect -407 5 -404 13
rect -390 5 -387 13
rect -407 -9 -387 5
rect -407 -17 -404 -9
rect -390 -17 -387 -9
rect -63 -29 -57 -11
rect -29 -29 -23 -11
rect -63 -40 -23 -29
rect -63 -58 -57 -40
rect -29 -58 -23 -40
rect -63 -73 -23 -58
rect -63 -91 -57 -73
rect -29 -91 -23 -73
rect 27 -29 33 -11
rect 61 -29 67 -11
rect 27 -40 67 -29
rect 27 -58 33 -40
rect 61 -58 67 -40
rect 27 -73 67 -58
rect 27 -91 33 -73
rect 61 -91 67 -73
rect 197 -29 203 -11
rect 231 -29 237 -11
rect 197 -40 237 -29
rect 197 -58 203 -40
rect 231 -58 237 -40
rect 197 -73 237 -58
rect 197 -91 203 -73
rect 231 -91 237 -73
rect 287 -29 293 -11
rect 321 -29 327 -11
rect 287 -40 327 -29
rect 287 -58 293 -40
rect 321 -58 327 -40
rect 287 -73 327 -58
rect 287 -91 293 -73
rect 321 -91 327 -73
<< pdiffusion >>
rect -503 180 -497 198
rect -469 180 -463 198
rect -503 159 -463 180
rect -503 141 -497 159
rect -469 141 -463 159
rect -503 116 -463 141
rect -503 98 -497 116
rect -469 98 -463 116
rect -413 180 -407 198
rect -379 180 -373 198
rect -413 159 -373 180
rect -413 141 -407 159
rect -379 141 -373 159
rect -413 116 -373 141
rect -243 184 -241 198
rect -225 184 -223 198
rect -243 167 -223 184
rect -243 153 -241 167
rect -225 153 -223 167
rect -243 132 -223 153
rect -243 118 -241 132
rect -225 118 -223 132
rect -213 184 -211 198
rect -195 184 -193 198
rect -213 167 -193 184
rect -213 153 -211 167
rect -195 153 -193 167
rect -213 132 -193 153
rect -213 118 -211 132
rect -195 118 -193 132
rect -63 180 -57 198
rect -29 180 -23 198
rect -63 151 -23 180
rect -63 133 -57 151
rect -29 133 -23 151
rect -413 98 -407 116
rect -379 98 -373 116
rect -63 96 -23 133
rect -63 78 -57 96
rect -29 78 -23 96
rect 27 180 33 198
rect 61 180 67 198
rect 27 151 67 180
rect 27 133 33 151
rect 61 133 67 151
rect 27 96 67 133
rect 27 78 33 96
rect 61 78 67 96
rect 197 180 203 198
rect 231 180 237 198
rect 197 151 237 180
rect 197 133 203 151
rect 231 133 237 151
rect 197 96 237 133
rect 197 78 203 96
rect 231 78 237 96
rect 287 180 293 198
rect 321 180 327 198
rect 287 151 327 180
rect 287 133 293 151
rect 321 133 327 151
rect 287 96 327 133
rect 287 78 293 96
rect 321 78 327 96
rect 457 180 463 198
rect 491 180 497 198
rect 457 151 497 180
rect 457 133 463 151
rect 491 133 497 151
rect 457 96 497 133
rect 457 78 463 96
rect 491 78 497 96
rect 547 180 553 198
rect 581 180 587 198
rect 547 151 587 180
rect 547 133 553 151
rect 581 133 587 151
rect 547 96 587 133
rect 547 78 553 96
rect 581 78 587 96
<< ndcontact >>
rect -494 5 -480 13
rect -494 -17 -480 -9
rect -464 5 -450 13
rect -464 -17 -450 -9
rect -434 5 -420 13
rect -434 -17 -420 -9
rect -404 5 -390 13
rect -404 -17 -390 -9
rect -57 -29 -29 -11
rect -57 -58 -29 -40
rect -57 -91 -29 -73
rect 33 -29 61 -11
rect 33 -58 61 -40
rect 33 -91 61 -73
rect 203 -29 231 -11
rect 203 -58 231 -40
rect 203 -91 231 -73
rect 293 -29 321 -11
rect 293 -58 321 -40
rect 293 -91 321 -73
<< pdcontact >>
rect -497 180 -469 198
rect -497 141 -469 159
rect -497 98 -469 116
rect -407 180 -379 198
rect -407 141 -379 159
rect -241 184 -225 198
rect -241 153 -225 167
rect -241 118 -225 132
rect -211 184 -195 198
rect -211 153 -195 167
rect -211 118 -195 132
rect -57 180 -29 198
rect -57 133 -29 151
rect -407 98 -379 116
rect -57 78 -29 96
rect 33 180 61 198
rect 33 133 61 151
rect 33 78 61 96
rect 203 180 231 198
rect 203 133 231 151
rect 203 78 231 96
rect 293 180 321 198
rect 293 133 321 151
rect 293 78 321 96
rect 463 180 491 198
rect 463 133 491 151
rect 463 78 491 96
rect 553 180 581 198
rect 553 133 581 151
rect 553 78 581 96
<< nsubstratencontact >>
rect -523 278 -497 308
rect -451 278 -425 308
rect -383 278 -357 308
rect -260 278 -234 308
rect -202 278 -176 308
rect -80 278 -54 308
rect -6 278 20 308
rect 58 278 84 308
rect 180 278 206 308
rect 251 278 277 308
rect 318 278 344 308
rect 440 278 466 308
rect 510 278 536 308
rect 578 278 604 308
<< polysilicon >>
rect -449 229 -445 241
rect -431 229 -427 241
rect -463 198 -413 229
rect -12 229 -4 241
rect 7 229 16 241
rect -223 198 -213 201
rect -23 198 27 229
rect 248 229 257 241
rect 268 229 276 241
rect 237 198 287 229
rect 508 229 517 241
rect 528 229 535 241
rect 497 201 546 229
rect 497 198 547 201
rect -463 95 -413 98
rect -223 64 -213 118
rect -23 75 27 78
rect 237 68 287 78
rect 497 68 547 78
rect -477 19 -464 24
rect -447 19 -434 24
rect -417 19 -404 24
rect -477 13 -467 19
rect -447 13 -437 19
rect -417 13 -407 19
rect -9 13 -5 29
rect 9 13 13 29
rect -23 -11 27 13
rect 251 13 255 29
rect 269 13 273 29
rect 237 -11 287 13
rect -477 -20 -467 -17
rect -447 -20 -437 -17
rect -417 -20 -407 -17
rect -23 -94 27 -91
rect 237 -94 287 -91
<< polycontact >>
rect -463 229 -449 241
rect -445 229 -431 241
rect -427 229 -413 241
rect -23 229 -12 241
rect -4 229 7 241
rect 16 229 27 241
rect 237 229 248 241
rect 257 229 268 241
rect 276 229 287 241
rect 497 229 508 241
rect 517 229 528 241
rect 535 229 546 241
rect -233 64 -223 74
rect -464 19 -450 24
rect -434 19 -420 24
rect -404 19 -390 24
rect -23 13 -9 29
rect -5 13 9 29
rect 13 13 27 29
rect 237 13 251 29
rect 255 13 269 29
rect 273 13 287 29
<< metal1 >>
rect -497 278 -451 308
rect -425 278 -383 308
rect -357 278 -260 308
rect -234 278 -202 308
rect -176 278 -80 308
rect -54 278 -6 308
rect 20 278 58 308
rect 84 278 180 308
rect 206 278 251 308
rect 277 278 318 308
rect 344 278 440 308
rect 466 278 510 308
rect 536 278 578 308
rect 604 278 607 308
rect -497 198 -469 278
rect -449 229 -445 241
rect -431 229 -427 241
rect -413 229 -82 241
rect -241 198 -225 229
rect -57 198 -29 278
rect -12 229 -4 241
rect 7 229 16 241
rect 27 229 174 241
rect 203 198 231 278
rect 248 229 257 241
rect 268 229 276 241
rect 287 229 438 241
rect -497 159 -469 180
rect -497 116 -469 141
rect -407 159 -379 180
rect -407 116 -379 141
rect -241 167 -225 184
rect -241 132 -225 153
rect -211 167 -195 184
rect -211 132 -195 153
rect -404 74 -390 98
rect -404 64 -233 74
rect -404 24 -390 64
rect -464 13 -450 19
rect -494 -9 -480 5
rect -464 -9 -450 5
rect -434 13 -420 19
rect -434 -9 -420 5
rect -404 13 -390 19
rect -211 29 -195 118
rect -57 151 -29 180
rect -57 96 -29 133
rect 33 151 61 180
rect 33 96 61 133
rect 203 151 231 180
rect 203 96 231 133
rect 293 198 321 229
rect 293 151 321 180
rect 293 96 321 133
rect 463 198 491 278
rect 508 229 517 241
rect 528 229 535 241
rect 463 151 491 180
rect 463 96 491 133
rect 553 151 581 180
rect 553 96 581 133
rect 33 29 61 78
rect -211 13 -23 29
rect -9 13 -5 29
rect 9 13 13 29
rect 27 13 237 29
rect 251 13 255 29
rect 269 13 273 29
rect -404 -9 -390 5
rect 33 -11 61 13
rect 293 -11 321 78
rect -494 -43 -480 -17
rect -57 -40 -29 -29
rect -57 -73 -29 -58
rect 33 -40 61 -29
rect 33 -73 61 -58
rect 203 -40 231 -29
rect 203 -73 231 -58
rect 293 -40 321 -29
rect 293 -73 321 -58
rect -57 -178 -29 -91
rect 207 -106 227 -91
rect 558 -100 578 78
<< m2contact >>
rect -82 229 -71 241
rect -23 229 -12 241
rect 174 229 185 241
rect 237 229 248 241
rect 438 229 449 241
rect 497 229 508 241
<< metal2 >>
rect -71 229 -23 241
rect 185 229 237 241
rect 449 229 497 241
<< labels >>
rlabel metal1 -394 131 -394 131 1 a
rlabel metal1 -426 -1 -426 -1 1 b
rlabel metal1 -459 -2 -459 -2 1 c
rlabel ptransistor -438 153 -438 154 1 2
rlabel metal1 110 294 110 294 1 1
rlabel metal1 46 -65 46 -65 1 3
rlabel metal1 -43 -64 -43 -64 1 4
rlabel metal1 214 -65 214 -65 1 5
rlabel metal1 566 104 566 104 1 vref
rlabel metal1 -44 -131 -44 -131 1 4
<< end >>
