magic
tech scmos
timestamp 1594246348
<< ntransistor >>
rect -477 -17 -467 13
rect -447 -17 -437 13
rect -417 -17 -407 13
<< ndiffusion >>
rect -497 5 -494 13
rect -480 5 -477 13
rect -497 -9 -477 5
rect -497 -17 -494 -9
rect -480 -17 -477 -9
rect -467 5 -464 13
rect -450 5 -447 13
rect -467 -9 -447 5
rect -467 -17 -464 -9
rect -450 -17 -447 -9
rect -437 5 -434 13
rect -420 5 -417 13
rect -437 -9 -417 5
rect -437 -17 -434 -9
rect -420 -17 -417 -9
rect -407 5 -404 13
rect -390 5 -387 13
rect -407 -9 -387 5
rect -407 -17 -404 -9
rect -390 -17 -387 -9
<< ndcontact >>
rect -494 5 -480 13
rect -494 -17 -480 -9
rect -464 5 -450 13
rect -464 -17 -450 -9
rect -434 5 -420 13
rect -434 -17 -420 -9
rect -404 5 -390 13
rect -404 -17 -390 -9
<< polysilicon >>
rect -477 19 -464 24
rect -447 19 -434 24
rect -417 19 -404 24
rect -477 13 -467 19
rect -447 13 -437 19
rect -417 13 -407 19
rect -477 -20 -467 -17
rect -447 -20 -437 -17
rect -417 -20 -407 -17
<< polycontact >>
rect -464 19 -450 24
rect -434 19 -420 24
rect -404 19 -390 24
<< metal1 >>
rect -404 24 -390 36
rect -464 13 -450 19
rect -494 -9 -480 5
rect -464 -9 -450 5
rect -434 13 -420 19
rect -434 -9 -420 5
rect -404 13 -390 19
rect -404 -9 -390 5
rect -494 -34 -480 -17
<< labels >>
rlabel metal1 -426 -1 -426 -1 1 b
rlabel metal1 -459 -2 -459 -2 1 c
<< end >>
