MACRO bandgap
  ORIGIN 0 0 ;
  FOREIGN bandgap 0 0 ;
  SIZE 31.972 BY 37.6 ;
  PIN 6
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 16.54 22.56 16.58 29.688 ;
      LAYER M2 ;
        RECT 7.324 18.716 17.956 18.748 ;
      LAYER M3 ;
        RECT 8.14 9.624 8.18 16.752 ;
      LAYER M3 ;
        RECT 7.82 22.644 7.86 30.444 ;
      LAYER M3 ;
        RECT 16.54 18.732 16.58 22.596 ;
      LAYER M2 ;
        RECT 16.544 18.716 16.576 18.748 ;
      LAYER M2 ;
        RECT 8.144 18.716 8.176 18.748 ;
      LAYER M3 ;
        RECT 8.14 16.716 8.18 18.732 ;
      LAYER M2 ;
        RECT 7.824 18.716 7.856 18.748 ;
      LAYER M3 ;
        RECT 7.82 18.732 7.86 22.68 ;
    END
  END 6
  PIN 4
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 0.364 20.648 26.996 20.68 ;
      LAYER M3 ;
        RECT 8.22 10.38 8.26 17.508 ;
      LAYER M3 ;
        RECT 17.34 9.708 17.38 17.508 ;
      LAYER M3 ;
        RECT 8.22 10.396 8.26 10.436 ;
      LAYER M4 ;
        RECT 8.24 10.396 17.36 10.436 ;
      LAYER M3 ;
        RECT 17.34 10.396 17.38 10.436 ;
      LAYER M3 ;
        RECT 7.9 22.728 7.94 29.856 ;
      LAYER M2 ;
        RECT 8.224 20.648 8.256 20.68 ;
      LAYER M3 ;
        RECT 8.22 17.472 8.26 20.664 ;
      LAYER M2 ;
        RECT 7.904 20.648 7.936 20.68 ;
      LAYER M3 ;
        RECT 7.9 20.664 7.94 22.764 ;
    END
  END 4
  PIN 9
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 6.508 9.392 6.58 9.424 ;
    END
  END 9
  PIN 8
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 5.164 9.392 5.236 9.424 ;
      LAYER M3 ;
        RECT 7.74 22.56 7.78 29.688 ;
      LAYER M2 ;
        RECT 5.2 9.392 6.4 9.424 ;
      LAYER M3 ;
        RECT 6.38 9.408 6.42 22.596 ;
      LAYER M4 ;
        RECT 6.4 22.576 7.76 22.616 ;
      LAYER M3 ;
        RECT 7.74 22.576 7.78 22.616 ;
    END
  END 8
  PIN 10
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 0.044 0.068 0.116 0.1 ;
    END
  END 10
  PIN 2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 12.46 1.056 12.5 8.184 ;
      LAYER M3 ;
        RECT 15.02 1.14 15.06 8.268 ;
      LAYER M3 ;
        RECT 18.38 0.384 18.42 8.268 ;
      LAYER M3 ;
        RECT 15.02 1.156 15.06 1.196 ;
      LAYER M4 ;
        RECT 15.04 1.156 18.4 1.196 ;
      LAYER M3 ;
        RECT 18.38 1.156 18.42 1.196 ;
      LAYER M3 ;
        RECT 12.46 1.24 12.5 1.28 ;
      LAYER M2 ;
        RECT 12.48 1.244 15.04 1.276 ;
      LAYER M3 ;
        RECT 15.02 1.24 15.06 1.28 ;
      LAYER M3 ;
        RECT 17.18 9.54 17.22 16.668 ;
      LAYER M3 ;
        RECT 18.38 8.232 18.42 9.576 ;
      LAYER M4 ;
        RECT 17.2 9.556 18.4 9.596 ;
      LAYER M3 ;
        RECT 17.18 9.556 17.22 9.596 ;
    END
  END 2
  PIN 5
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 18.46 0.468 18.5 7.596 ;
      LAYER M3 ;
        RECT 17.26 9.624 17.3 16.752 ;
      LAYER M3 ;
        RECT 18.46 7.56 18.5 9.66 ;
      LAYER M4 ;
        RECT 17.28 9.64 18.48 9.68 ;
      LAYER M3 ;
        RECT 17.26 9.64 17.3 9.68 ;
    END
  END 5
  PIN 3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 12.38 0.3 12.42 7.428 ;
      LAYER M3 ;
        RECT 8.06 9.54 8.1 16.668 ;
      LAYER M3 ;
        RECT 12.38 7.392 12.42 9.576 ;
      LAYER M4 ;
        RECT 8.08 9.556 12.4 9.596 ;
      LAYER M3 ;
        RECT 8.06 9.556 8.1 9.596 ;
    END
  END 3
  PIN 7
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 7.66 22.476 7.7 29.604 ;
    END
  END 7
  OBS 
  LAYER M2 ;
        RECT 15.556 30.98 17.884 31.012 ;
  LAYER M3 ;
        RECT 16.46 22.476 16.5 29.604 ;
  LAYER M2 ;
        RECT 0.116 21.992 27.244 22.024 ;
  LAYER M2 ;
        RECT 27.396 12.164 31.804 12.196 ;
  LAYER M2 ;
        RECT 27.396 24.68 31.804 24.712 ;
  LAYER M2 ;
        RECT 27.396 37.196 31.804 37.228 ;
  LAYER M3 ;
        RECT 29.42 25.164 29.46 35.82 ;
  LAYER M2 ;
        RECT 0.116 30.98 15.404 31.012 ;
  LAYER M2 ;
        RECT 16.464 30.98 16.496 31.012 ;
  LAYER M3 ;
        RECT 16.46 29.568 16.5 30.996 ;
  LAYER M3 ;
        RECT 16.46 22.008 16.5 22.512 ;
  LAYER M2 ;
        RECT 16.464 21.992 16.496 22.024 ;
  LAYER M2 ;
        RECT 27.2 21.992 27.44 22.024 ;
  LAYER M1 ;
        RECT 27.424 12.18 27.456 22.008 ;
  LAYER M2 ;
        RECT 27.424 12.164 27.456 12.196 ;
  LAYER M1 ;
        RECT 27.424 22.008 27.456 24.696 ;
  LAYER M2 ;
        RECT 27.424 24.68 27.456 24.712 ;
  LAYER M1 ;
        RECT 27.424 24.696 27.456 37.212 ;
  LAYER M2 ;
        RECT 27.424 37.196 27.456 37.228 ;
  LAYER M2 ;
        RECT 29.424 24.68 29.456 24.712 ;
  LAYER M3 ;
        RECT 29.42 24.696 29.46 25.2 ;
  LAYER M2 ;
        RECT 15.36 30.98 15.6 31.012 ;
  LAYER M2 ;
        RECT 16.444 30.98 16.516 31.012 ;
  LAYER M3 ;
        RECT 16.46 30.96 16.5 31.032 ;
  LAYER M2 ;
        RECT 16.444 21.992 16.516 22.024 ;
  LAYER M3 ;
        RECT 16.46 21.972 16.5 22.044 ;
  LAYER M2 ;
        RECT 16.444 30.98 16.516 31.012 ;
  LAYER M3 ;
        RECT 16.46 30.96 16.5 31.032 ;
  LAYER M1 ;
        RECT 27.424 12.144 27.456 12.216 ;
  LAYER M2 ;
        RECT 27.404 12.164 27.476 12.196 ;
  LAYER M1 ;
        RECT 27.424 21.972 27.456 22.044 ;
  LAYER M2 ;
        RECT 27.404 21.992 27.476 22.024 ;
  LAYER M2 ;
        RECT 16.444 21.992 16.516 22.024 ;
  LAYER M3 ;
        RECT 16.46 21.972 16.5 22.044 ;
  LAYER M2 ;
        RECT 16.444 30.98 16.516 31.012 ;
  LAYER M3 ;
        RECT 16.46 30.96 16.5 31.032 ;
  LAYER M1 ;
        RECT 27.424 12.144 27.456 12.216 ;
  LAYER M2 ;
        RECT 27.404 12.164 27.476 12.196 ;
  LAYER M1 ;
        RECT 27.424 21.972 27.456 22.044 ;
  LAYER M2 ;
        RECT 27.404 21.992 27.476 22.024 ;
  LAYER M1 ;
        RECT 27.424 24.66 27.456 24.732 ;
  LAYER M2 ;
        RECT 27.404 24.68 27.476 24.712 ;
  LAYER M2 ;
        RECT 16.444 21.992 16.516 22.024 ;
  LAYER M3 ;
        RECT 16.46 21.972 16.5 22.044 ;
  LAYER M2 ;
        RECT 16.444 30.98 16.516 31.012 ;
  LAYER M3 ;
        RECT 16.46 30.96 16.5 31.032 ;
  LAYER M1 ;
        RECT 27.424 12.144 27.456 12.216 ;
  LAYER M2 ;
        RECT 27.404 12.164 27.476 12.196 ;
  LAYER M1 ;
        RECT 27.424 21.972 27.456 22.044 ;
  LAYER M2 ;
        RECT 27.404 21.992 27.476 22.024 ;
  LAYER M1 ;
        RECT 27.424 24.66 27.456 24.732 ;
  LAYER M2 ;
        RECT 27.404 24.68 27.476 24.712 ;
  LAYER M1 ;
        RECT 27.424 37.176 27.456 37.248 ;
  LAYER M2 ;
        RECT 27.404 37.196 27.476 37.228 ;
  LAYER M2 ;
        RECT 16.444 21.992 16.516 22.024 ;
  LAYER M3 ;
        RECT 16.46 21.972 16.5 22.044 ;
  LAYER M2 ;
        RECT 16.444 30.98 16.516 31.012 ;
  LAYER M3 ;
        RECT 16.46 30.96 16.5 31.032 ;
  LAYER M1 ;
        RECT 27.424 12.144 27.456 12.216 ;
  LAYER M2 ;
        RECT 27.404 12.164 27.476 12.196 ;
  LAYER M1 ;
        RECT 27.424 21.972 27.456 22.044 ;
  LAYER M2 ;
        RECT 27.404 21.992 27.476 22.024 ;
  LAYER M1 ;
        RECT 27.424 24.66 27.456 24.732 ;
  LAYER M2 ;
        RECT 27.404 24.68 27.476 24.712 ;
  LAYER M1 ;
        RECT 27.424 37.176 27.456 37.248 ;
  LAYER M2 ;
        RECT 27.404 37.196 27.476 37.228 ;
  LAYER M2 ;
        RECT 16.444 21.992 16.516 22.024 ;
  LAYER M3 ;
        RECT 16.46 21.972 16.5 22.044 ;
  LAYER M2 ;
        RECT 16.444 30.98 16.516 31.012 ;
  LAYER M3 ;
        RECT 16.46 30.96 16.5 31.032 ;
  LAYER M2 ;
        RECT 29.404 24.68 29.476 24.712 ;
  LAYER M3 ;
        RECT 29.42 24.66 29.46 24.732 ;
  LAYER M1 ;
        RECT 27.424 12.144 27.456 12.216 ;
  LAYER M2 ;
        RECT 27.404 12.164 27.476 12.196 ;
  LAYER M1 ;
        RECT 27.424 21.972 27.456 22.044 ;
  LAYER M2 ;
        RECT 27.404 21.992 27.476 22.024 ;
  LAYER M1 ;
        RECT 27.424 24.66 27.456 24.732 ;
  LAYER M2 ;
        RECT 27.404 24.68 27.476 24.712 ;
  LAYER M1 ;
        RECT 27.424 37.176 27.456 37.248 ;
  LAYER M2 ;
        RECT 27.404 37.196 27.476 37.228 ;
  LAYER M2 ;
        RECT 16.444 21.992 16.516 22.024 ;
  LAYER M3 ;
        RECT 16.46 21.972 16.5 22.044 ;
  LAYER M2 ;
        RECT 16.444 30.98 16.516 31.012 ;
  LAYER M3 ;
        RECT 16.46 30.96 16.5 31.032 ;
  LAYER M2 ;
        RECT 29.404 24.68 29.476 24.712 ;
  LAYER M3 ;
        RECT 29.42 24.66 29.46 24.732 ;
  LAYER M1 ;
        RECT 27.424 12.144 27.456 12.216 ;
  LAYER M2 ;
        RECT 27.404 12.164 27.476 12.196 ;
  LAYER M1 ;
        RECT 27.424 21.972 27.456 22.044 ;
  LAYER M2 ;
        RECT 27.404 21.992 27.476 22.024 ;
  LAYER M1 ;
        RECT 27.424 24.66 27.456 24.732 ;
  LAYER M2 ;
        RECT 27.404 24.68 27.476 24.712 ;
  LAYER M1 ;
        RECT 27.424 37.176 27.456 37.248 ;
  LAYER M2 ;
        RECT 27.404 37.196 27.476 37.228 ;
  LAYER M2 ;
        RECT 16.444 21.992 16.516 22.024 ;
  LAYER M3 ;
        RECT 16.46 21.972 16.5 22.044 ;
  LAYER M2 ;
        RECT 16.444 30.98 16.516 31.012 ;
  LAYER M3 ;
        RECT 16.46 30.96 16.5 31.032 ;
  LAYER M2 ;
        RECT 29.404 24.68 29.476 24.712 ;
  LAYER M3 ;
        RECT 29.42 24.66 29.46 24.732 ;
  LAYER M3 ;
        RECT 16.62 23.316 16.66 30.444 ;
  LAYER M2 ;
        RECT 0.364 21.404 26.996 21.436 ;
  LAYER M2 ;
        RECT 0.284 20.564 27.076 20.596 ;
  LAYER M2 ;
        RECT 7.244 18.632 18.036 18.664 ;
  LAYER M2 ;
        RECT 7.264 20.564 7.296 20.596 ;
  LAYER M3 ;
        RECT 7.26 18.648 7.3 20.58 ;
  LAYER M2 ;
        RECT 7.264 18.632 7.296 18.664 ;
  LAYER M2 ;
        RECT 7.244 18.632 7.316 18.664 ;
  LAYER M3 ;
        RECT 7.26 18.612 7.3 18.684 ;
  LAYER M2 ;
        RECT 7.244 20.564 7.316 20.596 ;
  LAYER M3 ;
        RECT 7.26 20.544 7.3 20.616 ;
  LAYER M2 ;
        RECT 7.244 18.632 7.316 18.664 ;
  LAYER M3 ;
        RECT 7.26 18.612 7.3 18.684 ;
  LAYER M2 ;
        RECT 7.244 20.564 7.316 20.596 ;
  LAYER M3 ;
        RECT 7.26 20.544 7.3 20.616 ;
  LAYER M2 ;
        RECT 7.324 19.472 17.956 19.504 ;
  LAYER M3 ;
        RECT 29.5 0.216 29.54 11.628 ;
  LAYER M3 ;
        RECT 14.94 0.384 14.98 7.512 ;
  LAYER M2 ;
        RECT 17.92 19.472 24 19.504 ;
  LAYER M3 ;
        RECT 23.98 16.8 24.02 19.488 ;
  LAYER M4 ;
        RECT 24 16.78 29.52 16.82 ;
  LAYER M5 ;
        RECT 29.488 11.592 29.552 16.8 ;
  LAYER M4 ;
        RECT 29.45 11.572 29.59 11.612 ;
  LAYER M3 ;
        RECT 29.5 11.572 29.54 11.612 ;
  LAYER M3 ;
        RECT 29.5 0.988 29.54 1.028 ;
  LAYER M4 ;
        RECT 24.336 0.988 29.52 1.028 ;
  LAYER M5 ;
        RECT 24.304 0.958 24.368 1.058 ;
  LAYER M6 ;
        RECT 24.156 0.976 24.516 1.04 ;
  LAYER M7 ;
        RECT 24.304 0.828 24.368 1.188 ;
  LAYER M8 ;
        RECT 14.976 0.976 24.336 1.04 ;
  LAYER M7 ;
        RECT 14.944 0.828 15.008 1.188 ;
  LAYER M6 ;
        RECT 14.796 0.976 15.156 1.04 ;
  LAYER M5 ;
        RECT 14.944 0.958 15.008 1.058 ;
  LAYER M4 ;
        RECT 14.898 0.988 15.038 1.028 ;
  LAYER M3 ;
        RECT 14.94 0.988 14.98 1.028 ;
  LAYER M2 ;
        RECT 23.964 19.472 24.036 19.504 ;
  LAYER M3 ;
        RECT 23.98 19.452 24.02 19.524 ;
  LAYER M3 ;
        RECT 23.98 16.76 24.02 16.84 ;
  LAYER M4 ;
        RECT 23.96 16.78 24.04 16.82 ;
  LAYER M3 ;
        RECT 29.5 11.552 29.54 11.632 ;
  LAYER M4 ;
        RECT 29.48 11.572 29.56 11.612 ;
  LAYER M4 ;
        RECT 29.48 11.572 29.56 11.612 ;
  LAYER M5 ;
        RECT 29.488 11.552 29.552 11.632 ;
  LAYER M4 ;
        RECT 29.48 16.78 29.56 16.82 ;
  LAYER M5 ;
        RECT 29.488 16.76 29.552 16.84 ;
  LAYER M2 ;
        RECT 23.964 19.472 24.036 19.504 ;
  LAYER M3 ;
        RECT 23.98 19.452 24.02 19.524 ;
  LAYER M3 ;
        RECT 14.94 0.968 14.98 1.048 ;
  LAYER M4 ;
        RECT 14.92 0.988 15 1.028 ;
  LAYER M3 ;
        RECT 23.98 16.76 24.02 16.84 ;
  LAYER M4 ;
        RECT 23.96 16.78 24.04 16.82 ;
  LAYER M3 ;
        RECT 29.5 0.968 29.54 1.048 ;
  LAYER M4 ;
        RECT 29.48 0.988 29.56 1.028 ;
  LAYER M4 ;
        RECT 14.936 0.988 15.016 1.028 ;
  LAYER M5 ;
        RECT 14.944 0.968 15.008 1.048 ;
  LAYER M4 ;
        RECT 24.296 0.988 24.376 1.028 ;
  LAYER M5 ;
        RECT 24.304 0.968 24.368 1.048 ;
  LAYER M4 ;
        RECT 29.48 16.78 29.56 16.82 ;
  LAYER M5 ;
        RECT 29.488 16.76 29.552 16.84 ;
  LAYER M5 ;
        RECT 14.944 0.956 15.008 1.06 ;
  LAYER M6 ;
        RECT 14.924 0.976 15.028 1.04 ;
  LAYER M5 ;
        RECT 24.304 0.956 24.368 1.06 ;
  LAYER M6 ;
        RECT 24.284 0.976 24.388 1.04 ;
  LAYER M6 ;
        RECT 14.924 0.976 15.028 1.04 ;
  LAYER M7 ;
        RECT 14.944 0.956 15.008 1.06 ;
  LAYER M6 ;
        RECT 24.284 0.976 24.388 1.04 ;
  LAYER M7 ;
        RECT 24.304 0.956 24.368 1.06 ;
  LAYER M7 ;
        RECT 14.944 0.956 15.008 1.06 ;
  LAYER M8 ;
        RECT 14.924 0.976 15.028 1.04 ;
  LAYER M7 ;
        RECT 24.304 0.956 24.368 1.06 ;
  LAYER M8 ;
        RECT 24.284 0.976 24.388 1.04 ;
  LAYER M2 ;
        RECT 23.964 19.472 24.036 19.504 ;
  LAYER M3 ;
        RECT 23.98 19.452 24.02 19.524 ;
  LAYER M3 ;
        RECT 23.98 16.76 24.02 16.84 ;
  LAYER M4 ;
        RECT 23.96 16.78 24.04 16.82 ;
  LAYER M3 ;
        RECT 29.5 0.968 29.54 1.048 ;
  LAYER M4 ;
        RECT 29.48 0.988 29.56 1.028 ;
  LAYER M4 ;
        RECT 29.48 16.78 29.56 16.82 ;
  LAYER M5 ;
        RECT 29.488 16.76 29.552 16.84 ;
  LAYER M3 ;
        RECT 29.42 0.132 29.46 10.788 ;
  LAYER M3 ;
        RECT 29.5 12.732 29.54 24.144 ;
  LAYER M3 ;
        RECT 29.42 10.752 29.46 12.516 ;
  LAYER M2 ;
        RECT 29.38 12.5 29.58 12.532 ;
  LAYER M3 ;
        RECT 29.5 12.516 29.54 12.768 ;
  LAYER M2 ;
        RECT 29.404 12.5 29.476 12.532 ;
  LAYER M3 ;
        RECT 29.42 12.48 29.46 12.552 ;
  LAYER M2 ;
        RECT 29.484 12.5 29.556 12.532 ;
  LAYER M3 ;
        RECT 29.5 12.48 29.54 12.552 ;
  LAYER M3 ;
        RECT 29.42 12.648 29.46 23.304 ;
  LAYER M3 ;
        RECT 29.5 25.248 29.54 36.66 ;
  LAYER M3 ;
        RECT 29.42 23.268 29.46 24.528 ;
  LAYER M2 ;
        RECT 29.38 24.512 29.58 24.544 ;
  LAYER M3 ;
        RECT 29.5 24.528 29.54 25.284 ;
  LAYER M2 ;
        RECT 29.404 24.512 29.476 24.544 ;
  LAYER M3 ;
        RECT 29.42 24.492 29.46 24.564 ;
  LAYER M2 ;
        RECT 29.484 24.512 29.556 24.544 ;
  LAYER M3 ;
        RECT 29.5 24.492 29.54 24.564 ;
  LAYER M2 ;
        RECT 4.012 18.296 4.084 18.328 ;
  LAYER M3 ;
        RECT 17.42 9.792 17.46 16.92 ;
  LAYER M2 ;
        RECT 4.08 18.296 17.44 18.328 ;
  LAYER M3 ;
        RECT 17.42 16.884 17.46 18.312 ;
  LAYER M2 ;
        RECT 17.404 18.296 17.476 18.328 ;
  LAYER M3 ;
        RECT 17.42 18.276 17.46 18.348 ;
  LAYER M2 ;
        RECT 17.404 18.296 17.476 18.328 ;
  LAYER M3 ;
        RECT 17.42 18.276 17.46 18.348 ;
  LAYER M1 ;
        RECT 15.824 22.476 15.856 23.22 ;
  LAYER M1 ;
        RECT 15.824 23.316 15.856 23.556 ;
  LAYER M1 ;
        RECT 15.824 23.652 15.856 24.396 ;
  LAYER M1 ;
        RECT 15.824 24.492 15.856 24.732 ;
  LAYER M1 ;
        RECT 15.824 24.828 15.856 25.572 ;
  LAYER M1 ;
        RECT 15.824 25.668 15.856 25.908 ;
  LAYER M1 ;
        RECT 15.824 26.004 15.856 26.748 ;
  LAYER M1 ;
        RECT 15.824 26.844 15.856 27.084 ;
  LAYER M1 ;
        RECT 15.824 27.18 15.856 27.924 ;
  LAYER M1 ;
        RECT 15.824 28.02 15.856 28.26 ;
  LAYER M1 ;
        RECT 15.824 28.356 15.856 29.1 ;
  LAYER M1 ;
        RECT 15.824 29.196 15.856 29.436 ;
  LAYER M1 ;
        RECT 15.824 29.532 15.856 30.276 ;
  LAYER M1 ;
        RECT 15.824 30.372 15.856 30.612 ;
  LAYER M1 ;
        RECT 15.824 30.876 15.856 31.116 ;
  LAYER M1 ;
        RECT 15.744 22.476 15.776 23.22 ;
  LAYER M1 ;
        RECT 15.744 23.652 15.776 24.396 ;
  LAYER M1 ;
        RECT 15.744 24.828 15.776 25.572 ;
  LAYER M1 ;
        RECT 15.744 26.004 15.776 26.748 ;
  LAYER M1 ;
        RECT 15.744 27.18 15.776 27.924 ;
  LAYER M1 ;
        RECT 15.744 28.356 15.776 29.1 ;
  LAYER M1 ;
        RECT 15.744 29.532 15.776 30.276 ;
  LAYER M1 ;
        RECT 15.904 22.476 15.936 23.22 ;
  LAYER M1 ;
        RECT 15.904 23.652 15.936 24.396 ;
  LAYER M1 ;
        RECT 15.904 24.828 15.936 25.572 ;
  LAYER M1 ;
        RECT 15.904 26.004 15.936 26.748 ;
  LAYER M1 ;
        RECT 15.904 27.18 15.936 27.924 ;
  LAYER M1 ;
        RECT 15.904 28.356 15.936 29.1 ;
  LAYER M1 ;
        RECT 15.904 29.532 15.936 30.276 ;
  LAYER M1 ;
        RECT 15.984 22.476 16.016 23.22 ;
  LAYER M1 ;
        RECT 15.984 23.316 16.016 23.556 ;
  LAYER M1 ;
        RECT 15.984 23.652 16.016 24.396 ;
  LAYER M1 ;
        RECT 15.984 24.492 16.016 24.732 ;
  LAYER M1 ;
        RECT 15.984 24.828 16.016 25.572 ;
  LAYER M1 ;
        RECT 15.984 25.668 16.016 25.908 ;
  LAYER M1 ;
        RECT 15.984 26.004 16.016 26.748 ;
  LAYER M1 ;
        RECT 15.984 26.844 16.016 27.084 ;
  LAYER M1 ;
        RECT 15.984 27.18 16.016 27.924 ;
  LAYER M1 ;
        RECT 15.984 28.02 16.016 28.26 ;
  LAYER M1 ;
        RECT 15.984 28.356 16.016 29.1 ;
  LAYER M1 ;
        RECT 15.984 29.196 16.016 29.436 ;
  LAYER M1 ;
        RECT 15.984 29.532 16.016 30.276 ;
  LAYER M1 ;
        RECT 15.984 30.372 16.016 30.612 ;
  LAYER M1 ;
        RECT 15.984 30.876 16.016 31.116 ;
  LAYER M1 ;
        RECT 16.064 22.476 16.096 23.22 ;
  LAYER M1 ;
        RECT 16.064 23.652 16.096 24.396 ;
  LAYER M1 ;
        RECT 16.064 24.828 16.096 25.572 ;
  LAYER M1 ;
        RECT 16.064 26.004 16.096 26.748 ;
  LAYER M1 ;
        RECT 16.064 27.18 16.096 27.924 ;
  LAYER M1 ;
        RECT 16.064 28.356 16.096 29.1 ;
  LAYER M1 ;
        RECT 16.064 29.532 16.096 30.276 ;
  LAYER M1 ;
        RECT 16.144 22.476 16.176 23.22 ;
  LAYER M1 ;
        RECT 16.144 23.316 16.176 23.556 ;
  LAYER M1 ;
        RECT 16.144 23.652 16.176 24.396 ;
  LAYER M1 ;
        RECT 16.144 24.492 16.176 24.732 ;
  LAYER M1 ;
        RECT 16.144 24.828 16.176 25.572 ;
  LAYER M1 ;
        RECT 16.144 25.668 16.176 25.908 ;
  LAYER M1 ;
        RECT 16.144 26.004 16.176 26.748 ;
  LAYER M1 ;
        RECT 16.144 26.844 16.176 27.084 ;
  LAYER M1 ;
        RECT 16.144 27.18 16.176 27.924 ;
  LAYER M1 ;
        RECT 16.144 28.02 16.176 28.26 ;
  LAYER M1 ;
        RECT 16.144 28.356 16.176 29.1 ;
  LAYER M1 ;
        RECT 16.144 29.196 16.176 29.436 ;
  LAYER M1 ;
        RECT 16.144 29.532 16.176 30.276 ;
  LAYER M1 ;
        RECT 16.144 30.372 16.176 30.612 ;
  LAYER M1 ;
        RECT 16.144 30.876 16.176 31.116 ;
  LAYER M1 ;
        RECT 16.224 22.476 16.256 23.22 ;
  LAYER M1 ;
        RECT 16.224 23.652 16.256 24.396 ;
  LAYER M1 ;
        RECT 16.224 24.828 16.256 25.572 ;
  LAYER M1 ;
        RECT 16.224 26.004 16.256 26.748 ;
  LAYER M1 ;
        RECT 16.224 27.18 16.256 27.924 ;
  LAYER M1 ;
        RECT 16.224 28.356 16.256 29.1 ;
  LAYER M1 ;
        RECT 16.224 29.532 16.256 30.276 ;
  LAYER M1 ;
        RECT 16.304 22.476 16.336 23.22 ;
  LAYER M1 ;
        RECT 16.304 23.316 16.336 23.556 ;
  LAYER M1 ;
        RECT 16.304 23.652 16.336 24.396 ;
  LAYER M1 ;
        RECT 16.304 24.492 16.336 24.732 ;
  LAYER M1 ;
        RECT 16.304 24.828 16.336 25.572 ;
  LAYER M1 ;
        RECT 16.304 25.668 16.336 25.908 ;
  LAYER M1 ;
        RECT 16.304 26.004 16.336 26.748 ;
  LAYER M1 ;
        RECT 16.304 26.844 16.336 27.084 ;
  LAYER M1 ;
        RECT 16.304 27.18 16.336 27.924 ;
  LAYER M1 ;
        RECT 16.304 28.02 16.336 28.26 ;
  LAYER M1 ;
        RECT 16.304 28.356 16.336 29.1 ;
  LAYER M1 ;
        RECT 16.304 29.196 16.336 29.436 ;
  LAYER M1 ;
        RECT 16.304 29.532 16.336 30.276 ;
  LAYER M1 ;
        RECT 16.304 30.372 16.336 30.612 ;
  LAYER M1 ;
        RECT 16.304 30.876 16.336 31.116 ;
  LAYER M1 ;
        RECT 16.384 22.476 16.416 23.22 ;
  LAYER M1 ;
        RECT 16.384 23.652 16.416 24.396 ;
  LAYER M1 ;
        RECT 16.384 24.828 16.416 25.572 ;
  LAYER M1 ;
        RECT 16.384 26.004 16.416 26.748 ;
  LAYER M1 ;
        RECT 16.384 27.18 16.416 27.924 ;
  LAYER M1 ;
        RECT 16.384 28.356 16.416 29.1 ;
  LAYER M1 ;
        RECT 16.384 29.532 16.416 30.276 ;
  LAYER M1 ;
        RECT 16.464 22.476 16.496 23.22 ;
  LAYER M1 ;
        RECT 16.464 23.316 16.496 23.556 ;
  LAYER M1 ;
        RECT 16.464 23.652 16.496 24.396 ;
  LAYER M1 ;
        RECT 16.464 24.492 16.496 24.732 ;
  LAYER M1 ;
        RECT 16.464 24.828 16.496 25.572 ;
  LAYER M1 ;
        RECT 16.464 25.668 16.496 25.908 ;
  LAYER M1 ;
        RECT 16.464 26.004 16.496 26.748 ;
  LAYER M1 ;
        RECT 16.464 26.844 16.496 27.084 ;
  LAYER M1 ;
        RECT 16.464 27.18 16.496 27.924 ;
  LAYER M1 ;
        RECT 16.464 28.02 16.496 28.26 ;
  LAYER M1 ;
        RECT 16.464 28.356 16.496 29.1 ;
  LAYER M1 ;
        RECT 16.464 29.196 16.496 29.436 ;
  LAYER M1 ;
        RECT 16.464 29.532 16.496 30.276 ;
  LAYER M1 ;
        RECT 16.464 30.372 16.496 30.612 ;
  LAYER M1 ;
        RECT 16.464 30.876 16.496 31.116 ;
  LAYER M1 ;
        RECT 16.544 22.476 16.576 23.22 ;
  LAYER M1 ;
        RECT 16.544 23.652 16.576 24.396 ;
  LAYER M1 ;
        RECT 16.544 24.828 16.576 25.572 ;
  LAYER M1 ;
        RECT 16.544 26.004 16.576 26.748 ;
  LAYER M1 ;
        RECT 16.544 27.18 16.576 27.924 ;
  LAYER M1 ;
        RECT 16.544 28.356 16.576 29.1 ;
  LAYER M1 ;
        RECT 16.544 29.532 16.576 30.276 ;
  LAYER M1 ;
        RECT 16.624 22.476 16.656 23.22 ;
  LAYER M1 ;
        RECT 16.624 23.316 16.656 23.556 ;
  LAYER M1 ;
        RECT 16.624 23.652 16.656 24.396 ;
  LAYER M1 ;
        RECT 16.624 24.492 16.656 24.732 ;
  LAYER M1 ;
        RECT 16.624 24.828 16.656 25.572 ;
  LAYER M1 ;
        RECT 16.624 25.668 16.656 25.908 ;
  LAYER M1 ;
        RECT 16.624 26.004 16.656 26.748 ;
  LAYER M1 ;
        RECT 16.624 26.844 16.656 27.084 ;
  LAYER M1 ;
        RECT 16.624 27.18 16.656 27.924 ;
  LAYER M1 ;
        RECT 16.624 28.02 16.656 28.26 ;
  LAYER M1 ;
        RECT 16.624 28.356 16.656 29.1 ;
  LAYER M1 ;
        RECT 16.624 29.196 16.656 29.436 ;
  LAYER M1 ;
        RECT 16.624 29.532 16.656 30.276 ;
  LAYER M1 ;
        RECT 16.624 30.372 16.656 30.612 ;
  LAYER M1 ;
        RECT 16.624 30.876 16.656 31.116 ;
  LAYER M1 ;
        RECT 16.704 22.476 16.736 23.22 ;
  LAYER M1 ;
        RECT 16.704 23.652 16.736 24.396 ;
  LAYER M1 ;
        RECT 16.704 24.828 16.736 25.572 ;
  LAYER M1 ;
        RECT 16.704 26.004 16.736 26.748 ;
  LAYER M1 ;
        RECT 16.704 27.18 16.736 27.924 ;
  LAYER M1 ;
        RECT 16.704 28.356 16.736 29.1 ;
  LAYER M1 ;
        RECT 16.704 29.532 16.736 30.276 ;
  LAYER M1 ;
        RECT 16.784 22.476 16.816 23.22 ;
  LAYER M1 ;
        RECT 16.784 23.316 16.816 23.556 ;
  LAYER M1 ;
        RECT 16.784 23.652 16.816 24.396 ;
  LAYER M1 ;
        RECT 16.784 24.492 16.816 24.732 ;
  LAYER M1 ;
        RECT 16.784 24.828 16.816 25.572 ;
  LAYER M1 ;
        RECT 16.784 25.668 16.816 25.908 ;
  LAYER M1 ;
        RECT 16.784 26.004 16.816 26.748 ;
  LAYER M1 ;
        RECT 16.784 26.844 16.816 27.084 ;
  LAYER M1 ;
        RECT 16.784 27.18 16.816 27.924 ;
  LAYER M1 ;
        RECT 16.784 28.02 16.816 28.26 ;
  LAYER M1 ;
        RECT 16.784 28.356 16.816 29.1 ;
  LAYER M1 ;
        RECT 16.784 29.196 16.816 29.436 ;
  LAYER M1 ;
        RECT 16.784 29.532 16.816 30.276 ;
  LAYER M1 ;
        RECT 16.784 30.372 16.816 30.612 ;
  LAYER M1 ;
        RECT 16.784 30.876 16.816 31.116 ;
  LAYER M1 ;
        RECT 16.864 22.476 16.896 23.22 ;
  LAYER M1 ;
        RECT 16.864 23.652 16.896 24.396 ;
  LAYER M1 ;
        RECT 16.864 24.828 16.896 25.572 ;
  LAYER M1 ;
        RECT 16.864 26.004 16.896 26.748 ;
  LAYER M1 ;
        RECT 16.864 27.18 16.896 27.924 ;
  LAYER M1 ;
        RECT 16.864 28.356 16.896 29.1 ;
  LAYER M1 ;
        RECT 16.864 29.532 16.896 30.276 ;
  LAYER M1 ;
        RECT 16.944 22.476 16.976 23.22 ;
  LAYER M1 ;
        RECT 16.944 23.316 16.976 23.556 ;
  LAYER M1 ;
        RECT 16.944 23.652 16.976 24.396 ;
  LAYER M1 ;
        RECT 16.944 24.492 16.976 24.732 ;
  LAYER M1 ;
        RECT 16.944 24.828 16.976 25.572 ;
  LAYER M1 ;
        RECT 16.944 25.668 16.976 25.908 ;
  LAYER M1 ;
        RECT 16.944 26.004 16.976 26.748 ;
  LAYER M1 ;
        RECT 16.944 26.844 16.976 27.084 ;
  LAYER M1 ;
        RECT 16.944 27.18 16.976 27.924 ;
  LAYER M1 ;
        RECT 16.944 28.02 16.976 28.26 ;
  LAYER M1 ;
        RECT 16.944 28.356 16.976 29.1 ;
  LAYER M1 ;
        RECT 16.944 29.196 16.976 29.436 ;
  LAYER M1 ;
        RECT 16.944 29.532 16.976 30.276 ;
  LAYER M1 ;
        RECT 16.944 30.372 16.976 30.612 ;
  LAYER M1 ;
        RECT 16.944 30.876 16.976 31.116 ;
  LAYER M1 ;
        RECT 17.024 22.476 17.056 23.22 ;
  LAYER M1 ;
        RECT 17.024 23.652 17.056 24.396 ;
  LAYER M1 ;
        RECT 17.024 24.828 17.056 25.572 ;
  LAYER M1 ;
        RECT 17.024 26.004 17.056 26.748 ;
  LAYER M1 ;
        RECT 17.024 27.18 17.056 27.924 ;
  LAYER M1 ;
        RECT 17.024 28.356 17.056 29.1 ;
  LAYER M1 ;
        RECT 17.024 29.532 17.056 30.276 ;
  LAYER M1 ;
        RECT 17.104 22.476 17.136 23.22 ;
  LAYER M1 ;
        RECT 17.104 23.316 17.136 23.556 ;
  LAYER M1 ;
        RECT 17.104 23.652 17.136 24.396 ;
  LAYER M1 ;
        RECT 17.104 24.492 17.136 24.732 ;
  LAYER M1 ;
        RECT 17.104 24.828 17.136 25.572 ;
  LAYER M1 ;
        RECT 17.104 25.668 17.136 25.908 ;
  LAYER M1 ;
        RECT 17.104 26.004 17.136 26.748 ;
  LAYER M1 ;
        RECT 17.104 26.844 17.136 27.084 ;
  LAYER M1 ;
        RECT 17.104 27.18 17.136 27.924 ;
  LAYER M1 ;
        RECT 17.104 28.02 17.136 28.26 ;
  LAYER M1 ;
        RECT 17.104 28.356 17.136 29.1 ;
  LAYER M1 ;
        RECT 17.104 29.196 17.136 29.436 ;
  LAYER M1 ;
        RECT 17.104 29.532 17.136 30.276 ;
  LAYER M1 ;
        RECT 17.104 30.372 17.136 30.612 ;
  LAYER M1 ;
        RECT 17.104 30.876 17.136 31.116 ;
  LAYER M1 ;
        RECT 17.184 22.476 17.216 23.22 ;
  LAYER M1 ;
        RECT 17.184 23.652 17.216 24.396 ;
  LAYER M1 ;
        RECT 17.184 24.828 17.216 25.572 ;
  LAYER M1 ;
        RECT 17.184 26.004 17.216 26.748 ;
  LAYER M1 ;
        RECT 17.184 27.18 17.216 27.924 ;
  LAYER M1 ;
        RECT 17.184 28.356 17.216 29.1 ;
  LAYER M1 ;
        RECT 17.184 29.532 17.216 30.276 ;
  LAYER M1 ;
        RECT 17.264 22.476 17.296 23.22 ;
  LAYER M1 ;
        RECT 17.264 23.316 17.296 23.556 ;
  LAYER M1 ;
        RECT 17.264 23.652 17.296 24.396 ;
  LAYER M1 ;
        RECT 17.264 24.492 17.296 24.732 ;
  LAYER M1 ;
        RECT 17.264 24.828 17.296 25.572 ;
  LAYER M1 ;
        RECT 17.264 25.668 17.296 25.908 ;
  LAYER M1 ;
        RECT 17.264 26.004 17.296 26.748 ;
  LAYER M1 ;
        RECT 17.264 26.844 17.296 27.084 ;
  LAYER M1 ;
        RECT 17.264 27.18 17.296 27.924 ;
  LAYER M1 ;
        RECT 17.264 28.02 17.296 28.26 ;
  LAYER M1 ;
        RECT 17.264 28.356 17.296 29.1 ;
  LAYER M1 ;
        RECT 17.264 29.196 17.296 29.436 ;
  LAYER M1 ;
        RECT 17.264 29.532 17.296 30.276 ;
  LAYER M1 ;
        RECT 17.264 30.372 17.296 30.612 ;
  LAYER M1 ;
        RECT 17.264 30.876 17.296 31.116 ;
  LAYER M1 ;
        RECT 17.344 22.476 17.376 23.22 ;
  LAYER M1 ;
        RECT 17.344 23.652 17.376 24.396 ;
  LAYER M1 ;
        RECT 17.344 24.828 17.376 25.572 ;
  LAYER M1 ;
        RECT 17.344 26.004 17.376 26.748 ;
  LAYER M1 ;
        RECT 17.344 27.18 17.376 27.924 ;
  LAYER M1 ;
        RECT 17.344 28.356 17.376 29.1 ;
  LAYER M1 ;
        RECT 17.344 29.532 17.376 30.276 ;
  LAYER M1 ;
        RECT 17.424 22.476 17.456 23.22 ;
  LAYER M1 ;
        RECT 17.424 23.316 17.456 23.556 ;
  LAYER M1 ;
        RECT 17.424 23.652 17.456 24.396 ;
  LAYER M1 ;
        RECT 17.424 24.492 17.456 24.732 ;
  LAYER M1 ;
        RECT 17.424 24.828 17.456 25.572 ;
  LAYER M1 ;
        RECT 17.424 25.668 17.456 25.908 ;
  LAYER M1 ;
        RECT 17.424 26.004 17.456 26.748 ;
  LAYER M1 ;
        RECT 17.424 26.844 17.456 27.084 ;
  LAYER M1 ;
        RECT 17.424 27.18 17.456 27.924 ;
  LAYER M1 ;
        RECT 17.424 28.02 17.456 28.26 ;
  LAYER M1 ;
        RECT 17.424 28.356 17.456 29.1 ;
  LAYER M1 ;
        RECT 17.424 29.196 17.456 29.436 ;
  LAYER M1 ;
        RECT 17.424 29.532 17.456 30.276 ;
  LAYER M1 ;
        RECT 17.424 30.372 17.456 30.612 ;
  LAYER M1 ;
        RECT 17.424 30.876 17.456 31.116 ;
  LAYER M1 ;
        RECT 17.504 22.476 17.536 23.22 ;
  LAYER M1 ;
        RECT 17.504 23.652 17.536 24.396 ;
  LAYER M1 ;
        RECT 17.504 24.828 17.536 25.572 ;
  LAYER M1 ;
        RECT 17.504 26.004 17.536 26.748 ;
  LAYER M1 ;
        RECT 17.504 27.18 17.536 27.924 ;
  LAYER M1 ;
        RECT 17.504 28.356 17.536 29.1 ;
  LAYER M1 ;
        RECT 17.504 29.532 17.536 30.276 ;
  LAYER M1 ;
        RECT 17.584 22.476 17.616 23.22 ;
  LAYER M1 ;
        RECT 17.584 23.316 17.616 23.556 ;
  LAYER M1 ;
        RECT 17.584 23.652 17.616 24.396 ;
  LAYER M1 ;
        RECT 17.584 24.492 17.616 24.732 ;
  LAYER M1 ;
        RECT 17.584 24.828 17.616 25.572 ;
  LAYER M1 ;
        RECT 17.584 25.668 17.616 25.908 ;
  LAYER M1 ;
        RECT 17.584 26.004 17.616 26.748 ;
  LAYER M1 ;
        RECT 17.584 26.844 17.616 27.084 ;
  LAYER M1 ;
        RECT 17.584 27.18 17.616 27.924 ;
  LAYER M1 ;
        RECT 17.584 28.02 17.616 28.26 ;
  LAYER M1 ;
        RECT 17.584 28.356 17.616 29.1 ;
  LAYER M1 ;
        RECT 17.584 29.196 17.616 29.436 ;
  LAYER M1 ;
        RECT 17.584 29.532 17.616 30.276 ;
  LAYER M1 ;
        RECT 17.584 30.372 17.616 30.612 ;
  LAYER M1 ;
        RECT 17.584 30.876 17.616 31.116 ;
  LAYER M1 ;
        RECT 17.664 22.476 17.696 23.22 ;
  LAYER M1 ;
        RECT 17.664 23.652 17.696 24.396 ;
  LAYER M1 ;
        RECT 17.664 24.828 17.696 25.572 ;
  LAYER M1 ;
        RECT 17.664 26.004 17.696 26.748 ;
  LAYER M1 ;
        RECT 17.664 27.18 17.696 27.924 ;
  LAYER M1 ;
        RECT 17.664 28.356 17.696 29.1 ;
  LAYER M1 ;
        RECT 17.664 29.532 17.696 30.276 ;
  LAYER M2 ;
        RECT 15.724 22.496 17.716 22.528 ;
  LAYER M2 ;
        RECT 15.804 22.58 17.636 22.612 ;
  LAYER M2 ;
        RECT 15.804 23.336 17.636 23.368 ;
  LAYER M2 ;
        RECT 15.724 23.672 17.716 23.704 ;
  LAYER M2 ;
        RECT 15.804 23.756 17.636 23.788 ;
  LAYER M2 ;
        RECT 15.804 24.512 17.636 24.544 ;
  LAYER M2 ;
        RECT 15.724 24.848 17.716 24.88 ;
  LAYER M2 ;
        RECT 15.804 24.932 17.636 24.964 ;
  LAYER M2 ;
        RECT 15.804 25.688 17.636 25.72 ;
  LAYER M2 ;
        RECT 15.724 26.024 17.716 26.056 ;
  LAYER M2 ;
        RECT 15.804 26.108 17.636 26.14 ;
  LAYER M2 ;
        RECT 15.804 26.864 17.636 26.896 ;
  LAYER M2 ;
        RECT 15.724 27.2 17.716 27.232 ;
  LAYER M2 ;
        RECT 15.804 27.284 17.636 27.316 ;
  LAYER M2 ;
        RECT 15.804 28.04 17.636 28.072 ;
  LAYER M2 ;
        RECT 15.724 28.376 17.716 28.408 ;
  LAYER M2 ;
        RECT 15.804 28.46 17.636 28.492 ;
  LAYER M2 ;
        RECT 15.804 29.216 17.636 29.248 ;
  LAYER M2 ;
        RECT 15.724 29.552 17.716 29.584 ;
  LAYER M2 ;
        RECT 15.804 29.636 17.636 29.668 ;
  LAYER M2 ;
        RECT 15.804 30.392 17.636 30.424 ;
  LAYER M1 ;
        RECT 0.384 20.544 0.416 21.288 ;
  LAYER M1 ;
        RECT 0.384 21.384 0.416 21.624 ;
  LAYER M1 ;
        RECT 0.384 21.888 0.416 22.128 ;
  LAYER M1 ;
        RECT 0.304 20.544 0.336 21.288 ;
  LAYER M1 ;
        RECT 0.464 20.544 0.496 21.288 ;
  LAYER M1 ;
        RECT 0.544 20.544 0.576 21.288 ;
  LAYER M1 ;
        RECT 0.544 21.384 0.576 21.624 ;
  LAYER M1 ;
        RECT 0.544 21.888 0.576 22.128 ;
  LAYER M1 ;
        RECT 0.624 20.544 0.656 21.288 ;
  LAYER M1 ;
        RECT 0.704 20.544 0.736 21.288 ;
  LAYER M1 ;
        RECT 0.704 21.384 0.736 21.624 ;
  LAYER M1 ;
        RECT 0.704 21.888 0.736 22.128 ;
  LAYER M1 ;
        RECT 0.784 20.544 0.816 21.288 ;
  LAYER M1 ;
        RECT 0.864 20.544 0.896 21.288 ;
  LAYER M1 ;
        RECT 0.864 21.384 0.896 21.624 ;
  LAYER M1 ;
        RECT 0.864 21.888 0.896 22.128 ;
  LAYER M1 ;
        RECT 0.944 20.544 0.976 21.288 ;
  LAYER M1 ;
        RECT 1.024 20.544 1.056 21.288 ;
  LAYER M1 ;
        RECT 1.024 21.384 1.056 21.624 ;
  LAYER M1 ;
        RECT 1.024 21.888 1.056 22.128 ;
  LAYER M1 ;
        RECT 1.104 20.544 1.136 21.288 ;
  LAYER M1 ;
        RECT 1.184 20.544 1.216 21.288 ;
  LAYER M1 ;
        RECT 1.184 21.384 1.216 21.624 ;
  LAYER M1 ;
        RECT 1.184 21.888 1.216 22.128 ;
  LAYER M1 ;
        RECT 1.264 20.544 1.296 21.288 ;
  LAYER M1 ;
        RECT 1.344 20.544 1.376 21.288 ;
  LAYER M1 ;
        RECT 1.344 21.384 1.376 21.624 ;
  LAYER M1 ;
        RECT 1.344 21.888 1.376 22.128 ;
  LAYER M1 ;
        RECT 1.424 20.544 1.456 21.288 ;
  LAYER M1 ;
        RECT 1.504 20.544 1.536 21.288 ;
  LAYER M1 ;
        RECT 1.504 21.384 1.536 21.624 ;
  LAYER M1 ;
        RECT 1.504 21.888 1.536 22.128 ;
  LAYER M1 ;
        RECT 1.584 20.544 1.616 21.288 ;
  LAYER M1 ;
        RECT 1.664 20.544 1.696 21.288 ;
  LAYER M1 ;
        RECT 1.664 21.384 1.696 21.624 ;
  LAYER M1 ;
        RECT 1.664 21.888 1.696 22.128 ;
  LAYER M1 ;
        RECT 1.744 20.544 1.776 21.288 ;
  LAYER M1 ;
        RECT 1.824 20.544 1.856 21.288 ;
  LAYER M1 ;
        RECT 1.824 21.384 1.856 21.624 ;
  LAYER M1 ;
        RECT 1.824 21.888 1.856 22.128 ;
  LAYER M1 ;
        RECT 1.904 20.544 1.936 21.288 ;
  LAYER M1 ;
        RECT 1.984 20.544 2.016 21.288 ;
  LAYER M1 ;
        RECT 1.984 21.384 2.016 21.624 ;
  LAYER M1 ;
        RECT 1.984 21.888 2.016 22.128 ;
  LAYER M1 ;
        RECT 2.064 20.544 2.096 21.288 ;
  LAYER M1 ;
        RECT 2.144 20.544 2.176 21.288 ;
  LAYER M1 ;
        RECT 2.144 21.384 2.176 21.624 ;
  LAYER M1 ;
        RECT 2.144 21.888 2.176 22.128 ;
  LAYER M1 ;
        RECT 2.224 20.544 2.256 21.288 ;
  LAYER M1 ;
        RECT 2.304 20.544 2.336 21.288 ;
  LAYER M1 ;
        RECT 2.304 21.384 2.336 21.624 ;
  LAYER M1 ;
        RECT 2.304 21.888 2.336 22.128 ;
  LAYER M1 ;
        RECT 2.384 20.544 2.416 21.288 ;
  LAYER M1 ;
        RECT 2.464 20.544 2.496 21.288 ;
  LAYER M1 ;
        RECT 2.464 21.384 2.496 21.624 ;
  LAYER M1 ;
        RECT 2.464 21.888 2.496 22.128 ;
  LAYER M1 ;
        RECT 2.544 20.544 2.576 21.288 ;
  LAYER M1 ;
        RECT 2.624 20.544 2.656 21.288 ;
  LAYER M1 ;
        RECT 2.624 21.384 2.656 21.624 ;
  LAYER M1 ;
        RECT 2.624 21.888 2.656 22.128 ;
  LAYER M1 ;
        RECT 2.704 20.544 2.736 21.288 ;
  LAYER M1 ;
        RECT 2.784 20.544 2.816 21.288 ;
  LAYER M1 ;
        RECT 2.784 21.384 2.816 21.624 ;
  LAYER M1 ;
        RECT 2.784 21.888 2.816 22.128 ;
  LAYER M1 ;
        RECT 2.864 20.544 2.896 21.288 ;
  LAYER M1 ;
        RECT 2.944 20.544 2.976 21.288 ;
  LAYER M1 ;
        RECT 2.944 21.384 2.976 21.624 ;
  LAYER M1 ;
        RECT 2.944 21.888 2.976 22.128 ;
  LAYER M1 ;
        RECT 3.024 20.544 3.056 21.288 ;
  LAYER M1 ;
        RECT 3.104 20.544 3.136 21.288 ;
  LAYER M1 ;
        RECT 3.104 21.384 3.136 21.624 ;
  LAYER M1 ;
        RECT 3.104 21.888 3.136 22.128 ;
  LAYER M1 ;
        RECT 3.184 20.544 3.216 21.288 ;
  LAYER M1 ;
        RECT 3.264 20.544 3.296 21.288 ;
  LAYER M1 ;
        RECT 3.264 21.384 3.296 21.624 ;
  LAYER M1 ;
        RECT 3.264 21.888 3.296 22.128 ;
  LAYER M1 ;
        RECT 3.344 20.544 3.376 21.288 ;
  LAYER M1 ;
        RECT 3.424 20.544 3.456 21.288 ;
  LAYER M1 ;
        RECT 3.424 21.384 3.456 21.624 ;
  LAYER M1 ;
        RECT 3.424 21.888 3.456 22.128 ;
  LAYER M1 ;
        RECT 3.504 20.544 3.536 21.288 ;
  LAYER M1 ;
        RECT 3.584 20.544 3.616 21.288 ;
  LAYER M1 ;
        RECT 3.584 21.384 3.616 21.624 ;
  LAYER M1 ;
        RECT 3.584 21.888 3.616 22.128 ;
  LAYER M1 ;
        RECT 3.664 20.544 3.696 21.288 ;
  LAYER M1 ;
        RECT 3.744 20.544 3.776 21.288 ;
  LAYER M1 ;
        RECT 3.744 21.384 3.776 21.624 ;
  LAYER M1 ;
        RECT 3.744 21.888 3.776 22.128 ;
  LAYER M1 ;
        RECT 3.824 20.544 3.856 21.288 ;
  LAYER M1 ;
        RECT 3.904 20.544 3.936 21.288 ;
  LAYER M1 ;
        RECT 3.904 21.384 3.936 21.624 ;
  LAYER M1 ;
        RECT 3.904 21.888 3.936 22.128 ;
  LAYER M1 ;
        RECT 3.984 20.544 4.016 21.288 ;
  LAYER M1 ;
        RECT 4.064 20.544 4.096 21.288 ;
  LAYER M1 ;
        RECT 4.064 21.384 4.096 21.624 ;
  LAYER M1 ;
        RECT 4.064 21.888 4.096 22.128 ;
  LAYER M1 ;
        RECT 4.144 20.544 4.176 21.288 ;
  LAYER M1 ;
        RECT 4.224 20.544 4.256 21.288 ;
  LAYER M1 ;
        RECT 4.224 21.384 4.256 21.624 ;
  LAYER M1 ;
        RECT 4.224 21.888 4.256 22.128 ;
  LAYER M1 ;
        RECT 4.304 20.544 4.336 21.288 ;
  LAYER M1 ;
        RECT 4.384 20.544 4.416 21.288 ;
  LAYER M1 ;
        RECT 4.384 21.384 4.416 21.624 ;
  LAYER M1 ;
        RECT 4.384 21.888 4.416 22.128 ;
  LAYER M1 ;
        RECT 4.464 20.544 4.496 21.288 ;
  LAYER M1 ;
        RECT 4.544 20.544 4.576 21.288 ;
  LAYER M1 ;
        RECT 4.544 21.384 4.576 21.624 ;
  LAYER M1 ;
        RECT 4.544 21.888 4.576 22.128 ;
  LAYER M1 ;
        RECT 4.624 20.544 4.656 21.288 ;
  LAYER M1 ;
        RECT 4.704 20.544 4.736 21.288 ;
  LAYER M1 ;
        RECT 4.704 21.384 4.736 21.624 ;
  LAYER M1 ;
        RECT 4.704 21.888 4.736 22.128 ;
  LAYER M1 ;
        RECT 4.784 20.544 4.816 21.288 ;
  LAYER M1 ;
        RECT 4.864 20.544 4.896 21.288 ;
  LAYER M1 ;
        RECT 4.864 21.384 4.896 21.624 ;
  LAYER M1 ;
        RECT 4.864 21.888 4.896 22.128 ;
  LAYER M1 ;
        RECT 4.944 20.544 4.976 21.288 ;
  LAYER M1 ;
        RECT 5.024 20.544 5.056 21.288 ;
  LAYER M1 ;
        RECT 5.024 21.384 5.056 21.624 ;
  LAYER M1 ;
        RECT 5.024 21.888 5.056 22.128 ;
  LAYER M1 ;
        RECT 5.104 20.544 5.136 21.288 ;
  LAYER M1 ;
        RECT 5.184 20.544 5.216 21.288 ;
  LAYER M1 ;
        RECT 5.184 21.384 5.216 21.624 ;
  LAYER M1 ;
        RECT 5.184 21.888 5.216 22.128 ;
  LAYER M1 ;
        RECT 5.264 20.544 5.296 21.288 ;
  LAYER M1 ;
        RECT 5.344 20.544 5.376 21.288 ;
  LAYER M1 ;
        RECT 5.344 21.384 5.376 21.624 ;
  LAYER M1 ;
        RECT 5.344 21.888 5.376 22.128 ;
  LAYER M1 ;
        RECT 5.424 20.544 5.456 21.288 ;
  LAYER M1 ;
        RECT 5.504 20.544 5.536 21.288 ;
  LAYER M1 ;
        RECT 5.504 21.384 5.536 21.624 ;
  LAYER M1 ;
        RECT 5.504 21.888 5.536 22.128 ;
  LAYER M1 ;
        RECT 5.584 20.544 5.616 21.288 ;
  LAYER M1 ;
        RECT 5.664 20.544 5.696 21.288 ;
  LAYER M1 ;
        RECT 5.664 21.384 5.696 21.624 ;
  LAYER M1 ;
        RECT 5.664 21.888 5.696 22.128 ;
  LAYER M1 ;
        RECT 5.744 20.544 5.776 21.288 ;
  LAYER M1 ;
        RECT 5.824 20.544 5.856 21.288 ;
  LAYER M1 ;
        RECT 5.824 21.384 5.856 21.624 ;
  LAYER M1 ;
        RECT 5.824 21.888 5.856 22.128 ;
  LAYER M1 ;
        RECT 5.904 20.544 5.936 21.288 ;
  LAYER M1 ;
        RECT 5.984 20.544 6.016 21.288 ;
  LAYER M1 ;
        RECT 5.984 21.384 6.016 21.624 ;
  LAYER M1 ;
        RECT 5.984 21.888 6.016 22.128 ;
  LAYER M1 ;
        RECT 6.064 20.544 6.096 21.288 ;
  LAYER M1 ;
        RECT 6.144 20.544 6.176 21.288 ;
  LAYER M1 ;
        RECT 6.144 21.384 6.176 21.624 ;
  LAYER M1 ;
        RECT 6.144 21.888 6.176 22.128 ;
  LAYER M1 ;
        RECT 6.224 20.544 6.256 21.288 ;
  LAYER M1 ;
        RECT 6.304 20.544 6.336 21.288 ;
  LAYER M1 ;
        RECT 6.304 21.384 6.336 21.624 ;
  LAYER M1 ;
        RECT 6.304 21.888 6.336 22.128 ;
  LAYER M1 ;
        RECT 6.384 20.544 6.416 21.288 ;
  LAYER M1 ;
        RECT 6.464 20.544 6.496 21.288 ;
  LAYER M1 ;
        RECT 6.464 21.384 6.496 21.624 ;
  LAYER M1 ;
        RECT 6.464 21.888 6.496 22.128 ;
  LAYER M1 ;
        RECT 6.544 20.544 6.576 21.288 ;
  LAYER M1 ;
        RECT 6.624 20.544 6.656 21.288 ;
  LAYER M1 ;
        RECT 6.624 21.384 6.656 21.624 ;
  LAYER M1 ;
        RECT 6.624 21.888 6.656 22.128 ;
  LAYER M1 ;
        RECT 6.704 20.544 6.736 21.288 ;
  LAYER M1 ;
        RECT 6.784 20.544 6.816 21.288 ;
  LAYER M1 ;
        RECT 6.784 21.384 6.816 21.624 ;
  LAYER M1 ;
        RECT 6.784 21.888 6.816 22.128 ;
  LAYER M1 ;
        RECT 6.864 20.544 6.896 21.288 ;
  LAYER M1 ;
        RECT 6.944 20.544 6.976 21.288 ;
  LAYER M1 ;
        RECT 6.944 21.384 6.976 21.624 ;
  LAYER M1 ;
        RECT 6.944 21.888 6.976 22.128 ;
  LAYER M1 ;
        RECT 7.024 20.544 7.056 21.288 ;
  LAYER M1 ;
        RECT 7.104 20.544 7.136 21.288 ;
  LAYER M1 ;
        RECT 7.104 21.384 7.136 21.624 ;
  LAYER M1 ;
        RECT 7.104 21.888 7.136 22.128 ;
  LAYER M1 ;
        RECT 7.184 20.544 7.216 21.288 ;
  LAYER M1 ;
        RECT 7.264 20.544 7.296 21.288 ;
  LAYER M1 ;
        RECT 7.264 21.384 7.296 21.624 ;
  LAYER M1 ;
        RECT 7.264 21.888 7.296 22.128 ;
  LAYER M1 ;
        RECT 7.344 20.544 7.376 21.288 ;
  LAYER M1 ;
        RECT 7.424 20.544 7.456 21.288 ;
  LAYER M1 ;
        RECT 7.424 21.384 7.456 21.624 ;
  LAYER M1 ;
        RECT 7.424 21.888 7.456 22.128 ;
  LAYER M1 ;
        RECT 7.504 20.544 7.536 21.288 ;
  LAYER M1 ;
        RECT 7.584 20.544 7.616 21.288 ;
  LAYER M1 ;
        RECT 7.584 21.384 7.616 21.624 ;
  LAYER M1 ;
        RECT 7.584 21.888 7.616 22.128 ;
  LAYER M1 ;
        RECT 7.664 20.544 7.696 21.288 ;
  LAYER M1 ;
        RECT 7.744 20.544 7.776 21.288 ;
  LAYER M1 ;
        RECT 7.744 21.384 7.776 21.624 ;
  LAYER M1 ;
        RECT 7.744 21.888 7.776 22.128 ;
  LAYER M1 ;
        RECT 7.824 20.544 7.856 21.288 ;
  LAYER M1 ;
        RECT 7.904 20.544 7.936 21.288 ;
  LAYER M1 ;
        RECT 7.904 21.384 7.936 21.624 ;
  LAYER M1 ;
        RECT 7.904 21.888 7.936 22.128 ;
  LAYER M1 ;
        RECT 7.984 20.544 8.016 21.288 ;
  LAYER M1 ;
        RECT 8.064 20.544 8.096 21.288 ;
  LAYER M1 ;
        RECT 8.064 21.384 8.096 21.624 ;
  LAYER M1 ;
        RECT 8.064 21.888 8.096 22.128 ;
  LAYER M1 ;
        RECT 8.144 20.544 8.176 21.288 ;
  LAYER M1 ;
        RECT 8.224 20.544 8.256 21.288 ;
  LAYER M1 ;
        RECT 8.224 21.384 8.256 21.624 ;
  LAYER M1 ;
        RECT 8.224 21.888 8.256 22.128 ;
  LAYER M1 ;
        RECT 8.304 20.544 8.336 21.288 ;
  LAYER M1 ;
        RECT 8.384 20.544 8.416 21.288 ;
  LAYER M1 ;
        RECT 8.384 21.384 8.416 21.624 ;
  LAYER M1 ;
        RECT 8.384 21.888 8.416 22.128 ;
  LAYER M1 ;
        RECT 8.464 20.544 8.496 21.288 ;
  LAYER M1 ;
        RECT 8.544 20.544 8.576 21.288 ;
  LAYER M1 ;
        RECT 8.544 21.384 8.576 21.624 ;
  LAYER M1 ;
        RECT 8.544 21.888 8.576 22.128 ;
  LAYER M1 ;
        RECT 8.624 20.544 8.656 21.288 ;
  LAYER M1 ;
        RECT 8.704 20.544 8.736 21.288 ;
  LAYER M1 ;
        RECT 8.704 21.384 8.736 21.624 ;
  LAYER M1 ;
        RECT 8.704 21.888 8.736 22.128 ;
  LAYER M1 ;
        RECT 8.784 20.544 8.816 21.288 ;
  LAYER M1 ;
        RECT 8.864 20.544 8.896 21.288 ;
  LAYER M1 ;
        RECT 8.864 21.384 8.896 21.624 ;
  LAYER M1 ;
        RECT 8.864 21.888 8.896 22.128 ;
  LAYER M1 ;
        RECT 8.944 20.544 8.976 21.288 ;
  LAYER M1 ;
        RECT 9.024 20.544 9.056 21.288 ;
  LAYER M1 ;
        RECT 9.024 21.384 9.056 21.624 ;
  LAYER M1 ;
        RECT 9.024 21.888 9.056 22.128 ;
  LAYER M1 ;
        RECT 9.104 20.544 9.136 21.288 ;
  LAYER M1 ;
        RECT 9.184 20.544 9.216 21.288 ;
  LAYER M1 ;
        RECT 9.184 21.384 9.216 21.624 ;
  LAYER M1 ;
        RECT 9.184 21.888 9.216 22.128 ;
  LAYER M1 ;
        RECT 9.264 20.544 9.296 21.288 ;
  LAYER M1 ;
        RECT 9.344 20.544 9.376 21.288 ;
  LAYER M1 ;
        RECT 9.344 21.384 9.376 21.624 ;
  LAYER M1 ;
        RECT 9.344 21.888 9.376 22.128 ;
  LAYER M1 ;
        RECT 9.424 20.544 9.456 21.288 ;
  LAYER M1 ;
        RECT 9.504 20.544 9.536 21.288 ;
  LAYER M1 ;
        RECT 9.504 21.384 9.536 21.624 ;
  LAYER M1 ;
        RECT 9.504 21.888 9.536 22.128 ;
  LAYER M1 ;
        RECT 9.584 20.544 9.616 21.288 ;
  LAYER M1 ;
        RECT 9.664 20.544 9.696 21.288 ;
  LAYER M1 ;
        RECT 9.664 21.384 9.696 21.624 ;
  LAYER M1 ;
        RECT 9.664 21.888 9.696 22.128 ;
  LAYER M1 ;
        RECT 9.744 20.544 9.776 21.288 ;
  LAYER M1 ;
        RECT 9.824 20.544 9.856 21.288 ;
  LAYER M1 ;
        RECT 9.824 21.384 9.856 21.624 ;
  LAYER M1 ;
        RECT 9.824 21.888 9.856 22.128 ;
  LAYER M1 ;
        RECT 9.904 20.544 9.936 21.288 ;
  LAYER M1 ;
        RECT 9.984 20.544 10.016 21.288 ;
  LAYER M1 ;
        RECT 9.984 21.384 10.016 21.624 ;
  LAYER M1 ;
        RECT 9.984 21.888 10.016 22.128 ;
  LAYER M1 ;
        RECT 10.064 20.544 10.096 21.288 ;
  LAYER M1 ;
        RECT 10.144 20.544 10.176 21.288 ;
  LAYER M1 ;
        RECT 10.144 21.384 10.176 21.624 ;
  LAYER M1 ;
        RECT 10.144 21.888 10.176 22.128 ;
  LAYER M1 ;
        RECT 10.224 20.544 10.256 21.288 ;
  LAYER M1 ;
        RECT 10.304 20.544 10.336 21.288 ;
  LAYER M1 ;
        RECT 10.304 21.384 10.336 21.624 ;
  LAYER M1 ;
        RECT 10.304 21.888 10.336 22.128 ;
  LAYER M1 ;
        RECT 10.384 20.544 10.416 21.288 ;
  LAYER M1 ;
        RECT 10.464 20.544 10.496 21.288 ;
  LAYER M1 ;
        RECT 10.464 21.384 10.496 21.624 ;
  LAYER M1 ;
        RECT 10.464 21.888 10.496 22.128 ;
  LAYER M1 ;
        RECT 10.544 20.544 10.576 21.288 ;
  LAYER M1 ;
        RECT 10.624 20.544 10.656 21.288 ;
  LAYER M1 ;
        RECT 10.624 21.384 10.656 21.624 ;
  LAYER M1 ;
        RECT 10.624 21.888 10.656 22.128 ;
  LAYER M1 ;
        RECT 10.704 20.544 10.736 21.288 ;
  LAYER M1 ;
        RECT 10.784 20.544 10.816 21.288 ;
  LAYER M1 ;
        RECT 10.784 21.384 10.816 21.624 ;
  LAYER M1 ;
        RECT 10.784 21.888 10.816 22.128 ;
  LAYER M1 ;
        RECT 10.864 20.544 10.896 21.288 ;
  LAYER M1 ;
        RECT 10.944 20.544 10.976 21.288 ;
  LAYER M1 ;
        RECT 10.944 21.384 10.976 21.624 ;
  LAYER M1 ;
        RECT 10.944 21.888 10.976 22.128 ;
  LAYER M1 ;
        RECT 11.024 20.544 11.056 21.288 ;
  LAYER M1 ;
        RECT 11.104 20.544 11.136 21.288 ;
  LAYER M1 ;
        RECT 11.104 21.384 11.136 21.624 ;
  LAYER M1 ;
        RECT 11.104 21.888 11.136 22.128 ;
  LAYER M1 ;
        RECT 11.184 20.544 11.216 21.288 ;
  LAYER M1 ;
        RECT 11.264 20.544 11.296 21.288 ;
  LAYER M1 ;
        RECT 11.264 21.384 11.296 21.624 ;
  LAYER M1 ;
        RECT 11.264 21.888 11.296 22.128 ;
  LAYER M1 ;
        RECT 11.344 20.544 11.376 21.288 ;
  LAYER M1 ;
        RECT 11.424 20.544 11.456 21.288 ;
  LAYER M1 ;
        RECT 11.424 21.384 11.456 21.624 ;
  LAYER M1 ;
        RECT 11.424 21.888 11.456 22.128 ;
  LAYER M1 ;
        RECT 11.504 20.544 11.536 21.288 ;
  LAYER M1 ;
        RECT 11.584 20.544 11.616 21.288 ;
  LAYER M1 ;
        RECT 11.584 21.384 11.616 21.624 ;
  LAYER M1 ;
        RECT 11.584 21.888 11.616 22.128 ;
  LAYER M1 ;
        RECT 11.664 20.544 11.696 21.288 ;
  LAYER M1 ;
        RECT 11.744 20.544 11.776 21.288 ;
  LAYER M1 ;
        RECT 11.744 21.384 11.776 21.624 ;
  LAYER M1 ;
        RECT 11.744 21.888 11.776 22.128 ;
  LAYER M1 ;
        RECT 11.824 20.544 11.856 21.288 ;
  LAYER M1 ;
        RECT 11.904 20.544 11.936 21.288 ;
  LAYER M1 ;
        RECT 11.904 21.384 11.936 21.624 ;
  LAYER M1 ;
        RECT 11.904 21.888 11.936 22.128 ;
  LAYER M1 ;
        RECT 11.984 20.544 12.016 21.288 ;
  LAYER M1 ;
        RECT 12.064 20.544 12.096 21.288 ;
  LAYER M1 ;
        RECT 12.064 21.384 12.096 21.624 ;
  LAYER M1 ;
        RECT 12.064 21.888 12.096 22.128 ;
  LAYER M1 ;
        RECT 12.144 20.544 12.176 21.288 ;
  LAYER M1 ;
        RECT 12.224 20.544 12.256 21.288 ;
  LAYER M1 ;
        RECT 12.224 21.384 12.256 21.624 ;
  LAYER M1 ;
        RECT 12.224 21.888 12.256 22.128 ;
  LAYER M1 ;
        RECT 12.304 20.544 12.336 21.288 ;
  LAYER M1 ;
        RECT 12.384 20.544 12.416 21.288 ;
  LAYER M1 ;
        RECT 12.384 21.384 12.416 21.624 ;
  LAYER M1 ;
        RECT 12.384 21.888 12.416 22.128 ;
  LAYER M1 ;
        RECT 12.464 20.544 12.496 21.288 ;
  LAYER M1 ;
        RECT 12.544 20.544 12.576 21.288 ;
  LAYER M1 ;
        RECT 12.544 21.384 12.576 21.624 ;
  LAYER M1 ;
        RECT 12.544 21.888 12.576 22.128 ;
  LAYER M1 ;
        RECT 12.624 20.544 12.656 21.288 ;
  LAYER M1 ;
        RECT 12.704 20.544 12.736 21.288 ;
  LAYER M1 ;
        RECT 12.704 21.384 12.736 21.624 ;
  LAYER M1 ;
        RECT 12.704 21.888 12.736 22.128 ;
  LAYER M1 ;
        RECT 12.784 20.544 12.816 21.288 ;
  LAYER M1 ;
        RECT 12.864 20.544 12.896 21.288 ;
  LAYER M1 ;
        RECT 12.864 21.384 12.896 21.624 ;
  LAYER M1 ;
        RECT 12.864 21.888 12.896 22.128 ;
  LAYER M1 ;
        RECT 12.944 20.544 12.976 21.288 ;
  LAYER M1 ;
        RECT 13.024 20.544 13.056 21.288 ;
  LAYER M1 ;
        RECT 13.024 21.384 13.056 21.624 ;
  LAYER M1 ;
        RECT 13.024 21.888 13.056 22.128 ;
  LAYER M1 ;
        RECT 13.104 20.544 13.136 21.288 ;
  LAYER M1 ;
        RECT 13.184 20.544 13.216 21.288 ;
  LAYER M1 ;
        RECT 13.184 21.384 13.216 21.624 ;
  LAYER M1 ;
        RECT 13.184 21.888 13.216 22.128 ;
  LAYER M1 ;
        RECT 13.264 20.544 13.296 21.288 ;
  LAYER M1 ;
        RECT 13.344 20.544 13.376 21.288 ;
  LAYER M1 ;
        RECT 13.344 21.384 13.376 21.624 ;
  LAYER M1 ;
        RECT 13.344 21.888 13.376 22.128 ;
  LAYER M1 ;
        RECT 13.424 20.544 13.456 21.288 ;
  LAYER M1 ;
        RECT 13.504 20.544 13.536 21.288 ;
  LAYER M1 ;
        RECT 13.504 21.384 13.536 21.624 ;
  LAYER M1 ;
        RECT 13.504 21.888 13.536 22.128 ;
  LAYER M1 ;
        RECT 13.584 20.544 13.616 21.288 ;
  LAYER M1 ;
        RECT 13.664 20.544 13.696 21.288 ;
  LAYER M1 ;
        RECT 13.664 21.384 13.696 21.624 ;
  LAYER M1 ;
        RECT 13.664 21.888 13.696 22.128 ;
  LAYER M1 ;
        RECT 13.744 20.544 13.776 21.288 ;
  LAYER M1 ;
        RECT 13.824 20.544 13.856 21.288 ;
  LAYER M1 ;
        RECT 13.824 21.384 13.856 21.624 ;
  LAYER M1 ;
        RECT 13.824 21.888 13.856 22.128 ;
  LAYER M1 ;
        RECT 13.904 20.544 13.936 21.288 ;
  LAYER M1 ;
        RECT 13.984 20.544 14.016 21.288 ;
  LAYER M1 ;
        RECT 13.984 21.384 14.016 21.624 ;
  LAYER M1 ;
        RECT 13.984 21.888 14.016 22.128 ;
  LAYER M1 ;
        RECT 14.064 20.544 14.096 21.288 ;
  LAYER M1 ;
        RECT 14.144 20.544 14.176 21.288 ;
  LAYER M1 ;
        RECT 14.144 21.384 14.176 21.624 ;
  LAYER M1 ;
        RECT 14.144 21.888 14.176 22.128 ;
  LAYER M1 ;
        RECT 14.224 20.544 14.256 21.288 ;
  LAYER M1 ;
        RECT 14.304 20.544 14.336 21.288 ;
  LAYER M1 ;
        RECT 14.304 21.384 14.336 21.624 ;
  LAYER M1 ;
        RECT 14.304 21.888 14.336 22.128 ;
  LAYER M1 ;
        RECT 14.384 20.544 14.416 21.288 ;
  LAYER M1 ;
        RECT 14.464 20.544 14.496 21.288 ;
  LAYER M1 ;
        RECT 14.464 21.384 14.496 21.624 ;
  LAYER M1 ;
        RECT 14.464 21.888 14.496 22.128 ;
  LAYER M1 ;
        RECT 14.544 20.544 14.576 21.288 ;
  LAYER M1 ;
        RECT 14.624 20.544 14.656 21.288 ;
  LAYER M1 ;
        RECT 14.624 21.384 14.656 21.624 ;
  LAYER M1 ;
        RECT 14.624 21.888 14.656 22.128 ;
  LAYER M1 ;
        RECT 14.704 20.544 14.736 21.288 ;
  LAYER M1 ;
        RECT 14.784 20.544 14.816 21.288 ;
  LAYER M1 ;
        RECT 14.784 21.384 14.816 21.624 ;
  LAYER M1 ;
        RECT 14.784 21.888 14.816 22.128 ;
  LAYER M1 ;
        RECT 14.864 20.544 14.896 21.288 ;
  LAYER M1 ;
        RECT 14.944 20.544 14.976 21.288 ;
  LAYER M1 ;
        RECT 14.944 21.384 14.976 21.624 ;
  LAYER M1 ;
        RECT 14.944 21.888 14.976 22.128 ;
  LAYER M1 ;
        RECT 15.024 20.544 15.056 21.288 ;
  LAYER M1 ;
        RECT 15.104 20.544 15.136 21.288 ;
  LAYER M1 ;
        RECT 15.104 21.384 15.136 21.624 ;
  LAYER M1 ;
        RECT 15.104 21.888 15.136 22.128 ;
  LAYER M1 ;
        RECT 15.184 20.544 15.216 21.288 ;
  LAYER M1 ;
        RECT 15.264 20.544 15.296 21.288 ;
  LAYER M1 ;
        RECT 15.264 21.384 15.296 21.624 ;
  LAYER M1 ;
        RECT 15.264 21.888 15.296 22.128 ;
  LAYER M1 ;
        RECT 15.344 20.544 15.376 21.288 ;
  LAYER M1 ;
        RECT 15.424 20.544 15.456 21.288 ;
  LAYER M1 ;
        RECT 15.424 21.384 15.456 21.624 ;
  LAYER M1 ;
        RECT 15.424 21.888 15.456 22.128 ;
  LAYER M1 ;
        RECT 15.504 20.544 15.536 21.288 ;
  LAYER M1 ;
        RECT 15.584 20.544 15.616 21.288 ;
  LAYER M1 ;
        RECT 15.584 21.384 15.616 21.624 ;
  LAYER M1 ;
        RECT 15.584 21.888 15.616 22.128 ;
  LAYER M1 ;
        RECT 15.664 20.544 15.696 21.288 ;
  LAYER M1 ;
        RECT 15.744 20.544 15.776 21.288 ;
  LAYER M1 ;
        RECT 15.744 21.384 15.776 21.624 ;
  LAYER M1 ;
        RECT 15.744 21.888 15.776 22.128 ;
  LAYER M1 ;
        RECT 15.824 20.544 15.856 21.288 ;
  LAYER M1 ;
        RECT 15.904 20.544 15.936 21.288 ;
  LAYER M1 ;
        RECT 15.904 21.384 15.936 21.624 ;
  LAYER M1 ;
        RECT 15.904 21.888 15.936 22.128 ;
  LAYER M1 ;
        RECT 15.984 20.544 16.016 21.288 ;
  LAYER M1 ;
        RECT 16.064 20.544 16.096 21.288 ;
  LAYER M1 ;
        RECT 16.064 21.384 16.096 21.624 ;
  LAYER M1 ;
        RECT 16.064 21.888 16.096 22.128 ;
  LAYER M1 ;
        RECT 16.144 20.544 16.176 21.288 ;
  LAYER M1 ;
        RECT 16.224 20.544 16.256 21.288 ;
  LAYER M1 ;
        RECT 16.224 21.384 16.256 21.624 ;
  LAYER M1 ;
        RECT 16.224 21.888 16.256 22.128 ;
  LAYER M1 ;
        RECT 16.304 20.544 16.336 21.288 ;
  LAYER M1 ;
        RECT 16.384 20.544 16.416 21.288 ;
  LAYER M1 ;
        RECT 16.384 21.384 16.416 21.624 ;
  LAYER M1 ;
        RECT 16.384 21.888 16.416 22.128 ;
  LAYER M1 ;
        RECT 16.464 20.544 16.496 21.288 ;
  LAYER M1 ;
        RECT 16.544 20.544 16.576 21.288 ;
  LAYER M1 ;
        RECT 16.544 21.384 16.576 21.624 ;
  LAYER M1 ;
        RECT 16.544 21.888 16.576 22.128 ;
  LAYER M1 ;
        RECT 16.624 20.544 16.656 21.288 ;
  LAYER M1 ;
        RECT 16.704 20.544 16.736 21.288 ;
  LAYER M1 ;
        RECT 16.704 21.384 16.736 21.624 ;
  LAYER M1 ;
        RECT 16.704 21.888 16.736 22.128 ;
  LAYER M1 ;
        RECT 16.784 20.544 16.816 21.288 ;
  LAYER M1 ;
        RECT 16.864 20.544 16.896 21.288 ;
  LAYER M1 ;
        RECT 16.864 21.384 16.896 21.624 ;
  LAYER M1 ;
        RECT 16.864 21.888 16.896 22.128 ;
  LAYER M1 ;
        RECT 16.944 20.544 16.976 21.288 ;
  LAYER M1 ;
        RECT 17.024 20.544 17.056 21.288 ;
  LAYER M1 ;
        RECT 17.024 21.384 17.056 21.624 ;
  LAYER M1 ;
        RECT 17.024 21.888 17.056 22.128 ;
  LAYER M1 ;
        RECT 17.104 20.544 17.136 21.288 ;
  LAYER M1 ;
        RECT 17.184 20.544 17.216 21.288 ;
  LAYER M1 ;
        RECT 17.184 21.384 17.216 21.624 ;
  LAYER M1 ;
        RECT 17.184 21.888 17.216 22.128 ;
  LAYER M1 ;
        RECT 17.264 20.544 17.296 21.288 ;
  LAYER M1 ;
        RECT 17.344 20.544 17.376 21.288 ;
  LAYER M1 ;
        RECT 17.344 21.384 17.376 21.624 ;
  LAYER M1 ;
        RECT 17.344 21.888 17.376 22.128 ;
  LAYER M1 ;
        RECT 17.424 20.544 17.456 21.288 ;
  LAYER M1 ;
        RECT 17.504 20.544 17.536 21.288 ;
  LAYER M1 ;
        RECT 17.504 21.384 17.536 21.624 ;
  LAYER M1 ;
        RECT 17.504 21.888 17.536 22.128 ;
  LAYER M1 ;
        RECT 17.584 20.544 17.616 21.288 ;
  LAYER M1 ;
        RECT 17.664 20.544 17.696 21.288 ;
  LAYER M1 ;
        RECT 17.664 21.384 17.696 21.624 ;
  LAYER M1 ;
        RECT 17.664 21.888 17.696 22.128 ;
  LAYER M1 ;
        RECT 17.744 20.544 17.776 21.288 ;
  LAYER M1 ;
        RECT 17.824 20.544 17.856 21.288 ;
  LAYER M1 ;
        RECT 17.824 21.384 17.856 21.624 ;
  LAYER M1 ;
        RECT 17.824 21.888 17.856 22.128 ;
  LAYER M1 ;
        RECT 17.904 20.544 17.936 21.288 ;
  LAYER M1 ;
        RECT 17.984 20.544 18.016 21.288 ;
  LAYER M1 ;
        RECT 17.984 21.384 18.016 21.624 ;
  LAYER M1 ;
        RECT 17.984 21.888 18.016 22.128 ;
  LAYER M1 ;
        RECT 18.064 20.544 18.096 21.288 ;
  LAYER M1 ;
        RECT 18.144 20.544 18.176 21.288 ;
  LAYER M1 ;
        RECT 18.144 21.384 18.176 21.624 ;
  LAYER M1 ;
        RECT 18.144 21.888 18.176 22.128 ;
  LAYER M1 ;
        RECT 18.224 20.544 18.256 21.288 ;
  LAYER M1 ;
        RECT 18.304 20.544 18.336 21.288 ;
  LAYER M1 ;
        RECT 18.304 21.384 18.336 21.624 ;
  LAYER M1 ;
        RECT 18.304 21.888 18.336 22.128 ;
  LAYER M1 ;
        RECT 18.384 20.544 18.416 21.288 ;
  LAYER M1 ;
        RECT 18.464 20.544 18.496 21.288 ;
  LAYER M1 ;
        RECT 18.464 21.384 18.496 21.624 ;
  LAYER M1 ;
        RECT 18.464 21.888 18.496 22.128 ;
  LAYER M1 ;
        RECT 18.544 20.544 18.576 21.288 ;
  LAYER M1 ;
        RECT 18.624 20.544 18.656 21.288 ;
  LAYER M1 ;
        RECT 18.624 21.384 18.656 21.624 ;
  LAYER M1 ;
        RECT 18.624 21.888 18.656 22.128 ;
  LAYER M1 ;
        RECT 18.704 20.544 18.736 21.288 ;
  LAYER M1 ;
        RECT 18.784 20.544 18.816 21.288 ;
  LAYER M1 ;
        RECT 18.784 21.384 18.816 21.624 ;
  LAYER M1 ;
        RECT 18.784 21.888 18.816 22.128 ;
  LAYER M1 ;
        RECT 18.864 20.544 18.896 21.288 ;
  LAYER M1 ;
        RECT 18.944 20.544 18.976 21.288 ;
  LAYER M1 ;
        RECT 18.944 21.384 18.976 21.624 ;
  LAYER M1 ;
        RECT 18.944 21.888 18.976 22.128 ;
  LAYER M1 ;
        RECT 19.024 20.544 19.056 21.288 ;
  LAYER M1 ;
        RECT 19.104 20.544 19.136 21.288 ;
  LAYER M1 ;
        RECT 19.104 21.384 19.136 21.624 ;
  LAYER M1 ;
        RECT 19.104 21.888 19.136 22.128 ;
  LAYER M1 ;
        RECT 19.184 20.544 19.216 21.288 ;
  LAYER M1 ;
        RECT 19.264 20.544 19.296 21.288 ;
  LAYER M1 ;
        RECT 19.264 21.384 19.296 21.624 ;
  LAYER M1 ;
        RECT 19.264 21.888 19.296 22.128 ;
  LAYER M1 ;
        RECT 19.344 20.544 19.376 21.288 ;
  LAYER M1 ;
        RECT 19.424 20.544 19.456 21.288 ;
  LAYER M1 ;
        RECT 19.424 21.384 19.456 21.624 ;
  LAYER M1 ;
        RECT 19.424 21.888 19.456 22.128 ;
  LAYER M1 ;
        RECT 19.504 20.544 19.536 21.288 ;
  LAYER M1 ;
        RECT 19.584 20.544 19.616 21.288 ;
  LAYER M1 ;
        RECT 19.584 21.384 19.616 21.624 ;
  LAYER M1 ;
        RECT 19.584 21.888 19.616 22.128 ;
  LAYER M1 ;
        RECT 19.664 20.544 19.696 21.288 ;
  LAYER M1 ;
        RECT 19.744 20.544 19.776 21.288 ;
  LAYER M1 ;
        RECT 19.744 21.384 19.776 21.624 ;
  LAYER M1 ;
        RECT 19.744 21.888 19.776 22.128 ;
  LAYER M1 ;
        RECT 19.824 20.544 19.856 21.288 ;
  LAYER M1 ;
        RECT 19.904 20.544 19.936 21.288 ;
  LAYER M1 ;
        RECT 19.904 21.384 19.936 21.624 ;
  LAYER M1 ;
        RECT 19.904 21.888 19.936 22.128 ;
  LAYER M1 ;
        RECT 19.984 20.544 20.016 21.288 ;
  LAYER M1 ;
        RECT 20.064 20.544 20.096 21.288 ;
  LAYER M1 ;
        RECT 20.064 21.384 20.096 21.624 ;
  LAYER M1 ;
        RECT 20.064 21.888 20.096 22.128 ;
  LAYER M1 ;
        RECT 20.144 20.544 20.176 21.288 ;
  LAYER M1 ;
        RECT 20.224 20.544 20.256 21.288 ;
  LAYER M1 ;
        RECT 20.224 21.384 20.256 21.624 ;
  LAYER M1 ;
        RECT 20.224 21.888 20.256 22.128 ;
  LAYER M1 ;
        RECT 20.304 20.544 20.336 21.288 ;
  LAYER M1 ;
        RECT 20.384 20.544 20.416 21.288 ;
  LAYER M1 ;
        RECT 20.384 21.384 20.416 21.624 ;
  LAYER M1 ;
        RECT 20.384 21.888 20.416 22.128 ;
  LAYER M1 ;
        RECT 20.464 20.544 20.496 21.288 ;
  LAYER M1 ;
        RECT 20.544 20.544 20.576 21.288 ;
  LAYER M1 ;
        RECT 20.544 21.384 20.576 21.624 ;
  LAYER M1 ;
        RECT 20.544 21.888 20.576 22.128 ;
  LAYER M1 ;
        RECT 20.624 20.544 20.656 21.288 ;
  LAYER M1 ;
        RECT 20.704 20.544 20.736 21.288 ;
  LAYER M1 ;
        RECT 20.704 21.384 20.736 21.624 ;
  LAYER M1 ;
        RECT 20.704 21.888 20.736 22.128 ;
  LAYER M1 ;
        RECT 20.784 20.544 20.816 21.288 ;
  LAYER M1 ;
        RECT 20.864 20.544 20.896 21.288 ;
  LAYER M1 ;
        RECT 20.864 21.384 20.896 21.624 ;
  LAYER M1 ;
        RECT 20.864 21.888 20.896 22.128 ;
  LAYER M1 ;
        RECT 20.944 20.544 20.976 21.288 ;
  LAYER M1 ;
        RECT 21.024 20.544 21.056 21.288 ;
  LAYER M1 ;
        RECT 21.024 21.384 21.056 21.624 ;
  LAYER M1 ;
        RECT 21.024 21.888 21.056 22.128 ;
  LAYER M1 ;
        RECT 21.104 20.544 21.136 21.288 ;
  LAYER M1 ;
        RECT 21.184 20.544 21.216 21.288 ;
  LAYER M1 ;
        RECT 21.184 21.384 21.216 21.624 ;
  LAYER M1 ;
        RECT 21.184 21.888 21.216 22.128 ;
  LAYER M1 ;
        RECT 21.264 20.544 21.296 21.288 ;
  LAYER M1 ;
        RECT 21.344 20.544 21.376 21.288 ;
  LAYER M1 ;
        RECT 21.344 21.384 21.376 21.624 ;
  LAYER M1 ;
        RECT 21.344 21.888 21.376 22.128 ;
  LAYER M1 ;
        RECT 21.424 20.544 21.456 21.288 ;
  LAYER M1 ;
        RECT 21.504 20.544 21.536 21.288 ;
  LAYER M1 ;
        RECT 21.504 21.384 21.536 21.624 ;
  LAYER M1 ;
        RECT 21.504 21.888 21.536 22.128 ;
  LAYER M1 ;
        RECT 21.584 20.544 21.616 21.288 ;
  LAYER M1 ;
        RECT 21.664 20.544 21.696 21.288 ;
  LAYER M1 ;
        RECT 21.664 21.384 21.696 21.624 ;
  LAYER M1 ;
        RECT 21.664 21.888 21.696 22.128 ;
  LAYER M1 ;
        RECT 21.744 20.544 21.776 21.288 ;
  LAYER M1 ;
        RECT 21.824 20.544 21.856 21.288 ;
  LAYER M1 ;
        RECT 21.824 21.384 21.856 21.624 ;
  LAYER M1 ;
        RECT 21.824 21.888 21.856 22.128 ;
  LAYER M1 ;
        RECT 21.904 20.544 21.936 21.288 ;
  LAYER M1 ;
        RECT 21.984 20.544 22.016 21.288 ;
  LAYER M1 ;
        RECT 21.984 21.384 22.016 21.624 ;
  LAYER M1 ;
        RECT 21.984 21.888 22.016 22.128 ;
  LAYER M1 ;
        RECT 22.064 20.544 22.096 21.288 ;
  LAYER M1 ;
        RECT 22.144 20.544 22.176 21.288 ;
  LAYER M1 ;
        RECT 22.144 21.384 22.176 21.624 ;
  LAYER M1 ;
        RECT 22.144 21.888 22.176 22.128 ;
  LAYER M1 ;
        RECT 22.224 20.544 22.256 21.288 ;
  LAYER M1 ;
        RECT 22.304 20.544 22.336 21.288 ;
  LAYER M1 ;
        RECT 22.304 21.384 22.336 21.624 ;
  LAYER M1 ;
        RECT 22.304 21.888 22.336 22.128 ;
  LAYER M1 ;
        RECT 22.384 20.544 22.416 21.288 ;
  LAYER M1 ;
        RECT 22.464 20.544 22.496 21.288 ;
  LAYER M1 ;
        RECT 22.464 21.384 22.496 21.624 ;
  LAYER M1 ;
        RECT 22.464 21.888 22.496 22.128 ;
  LAYER M1 ;
        RECT 22.544 20.544 22.576 21.288 ;
  LAYER M1 ;
        RECT 22.624 20.544 22.656 21.288 ;
  LAYER M1 ;
        RECT 22.624 21.384 22.656 21.624 ;
  LAYER M1 ;
        RECT 22.624 21.888 22.656 22.128 ;
  LAYER M1 ;
        RECT 22.704 20.544 22.736 21.288 ;
  LAYER M1 ;
        RECT 22.784 20.544 22.816 21.288 ;
  LAYER M1 ;
        RECT 22.784 21.384 22.816 21.624 ;
  LAYER M1 ;
        RECT 22.784 21.888 22.816 22.128 ;
  LAYER M1 ;
        RECT 22.864 20.544 22.896 21.288 ;
  LAYER M1 ;
        RECT 22.944 20.544 22.976 21.288 ;
  LAYER M1 ;
        RECT 22.944 21.384 22.976 21.624 ;
  LAYER M1 ;
        RECT 22.944 21.888 22.976 22.128 ;
  LAYER M1 ;
        RECT 23.024 20.544 23.056 21.288 ;
  LAYER M1 ;
        RECT 23.104 20.544 23.136 21.288 ;
  LAYER M1 ;
        RECT 23.104 21.384 23.136 21.624 ;
  LAYER M1 ;
        RECT 23.104 21.888 23.136 22.128 ;
  LAYER M1 ;
        RECT 23.184 20.544 23.216 21.288 ;
  LAYER M1 ;
        RECT 23.264 20.544 23.296 21.288 ;
  LAYER M1 ;
        RECT 23.264 21.384 23.296 21.624 ;
  LAYER M1 ;
        RECT 23.264 21.888 23.296 22.128 ;
  LAYER M1 ;
        RECT 23.344 20.544 23.376 21.288 ;
  LAYER M1 ;
        RECT 23.424 20.544 23.456 21.288 ;
  LAYER M1 ;
        RECT 23.424 21.384 23.456 21.624 ;
  LAYER M1 ;
        RECT 23.424 21.888 23.456 22.128 ;
  LAYER M1 ;
        RECT 23.504 20.544 23.536 21.288 ;
  LAYER M1 ;
        RECT 23.584 20.544 23.616 21.288 ;
  LAYER M1 ;
        RECT 23.584 21.384 23.616 21.624 ;
  LAYER M1 ;
        RECT 23.584 21.888 23.616 22.128 ;
  LAYER M1 ;
        RECT 23.664 20.544 23.696 21.288 ;
  LAYER M1 ;
        RECT 23.744 20.544 23.776 21.288 ;
  LAYER M1 ;
        RECT 23.744 21.384 23.776 21.624 ;
  LAYER M1 ;
        RECT 23.744 21.888 23.776 22.128 ;
  LAYER M1 ;
        RECT 23.824 20.544 23.856 21.288 ;
  LAYER M1 ;
        RECT 23.904 20.544 23.936 21.288 ;
  LAYER M1 ;
        RECT 23.904 21.384 23.936 21.624 ;
  LAYER M1 ;
        RECT 23.904 21.888 23.936 22.128 ;
  LAYER M1 ;
        RECT 23.984 20.544 24.016 21.288 ;
  LAYER M1 ;
        RECT 24.064 20.544 24.096 21.288 ;
  LAYER M1 ;
        RECT 24.064 21.384 24.096 21.624 ;
  LAYER M1 ;
        RECT 24.064 21.888 24.096 22.128 ;
  LAYER M1 ;
        RECT 24.144 20.544 24.176 21.288 ;
  LAYER M1 ;
        RECT 24.224 20.544 24.256 21.288 ;
  LAYER M1 ;
        RECT 24.224 21.384 24.256 21.624 ;
  LAYER M1 ;
        RECT 24.224 21.888 24.256 22.128 ;
  LAYER M1 ;
        RECT 24.304 20.544 24.336 21.288 ;
  LAYER M1 ;
        RECT 24.384 20.544 24.416 21.288 ;
  LAYER M1 ;
        RECT 24.384 21.384 24.416 21.624 ;
  LAYER M1 ;
        RECT 24.384 21.888 24.416 22.128 ;
  LAYER M1 ;
        RECT 24.464 20.544 24.496 21.288 ;
  LAYER M1 ;
        RECT 24.544 20.544 24.576 21.288 ;
  LAYER M1 ;
        RECT 24.544 21.384 24.576 21.624 ;
  LAYER M1 ;
        RECT 24.544 21.888 24.576 22.128 ;
  LAYER M1 ;
        RECT 24.624 20.544 24.656 21.288 ;
  LAYER M1 ;
        RECT 24.704 20.544 24.736 21.288 ;
  LAYER M1 ;
        RECT 24.704 21.384 24.736 21.624 ;
  LAYER M1 ;
        RECT 24.704 21.888 24.736 22.128 ;
  LAYER M1 ;
        RECT 24.784 20.544 24.816 21.288 ;
  LAYER M1 ;
        RECT 24.864 20.544 24.896 21.288 ;
  LAYER M1 ;
        RECT 24.864 21.384 24.896 21.624 ;
  LAYER M1 ;
        RECT 24.864 21.888 24.896 22.128 ;
  LAYER M1 ;
        RECT 24.944 20.544 24.976 21.288 ;
  LAYER M1 ;
        RECT 25.024 20.544 25.056 21.288 ;
  LAYER M1 ;
        RECT 25.024 21.384 25.056 21.624 ;
  LAYER M1 ;
        RECT 25.024 21.888 25.056 22.128 ;
  LAYER M1 ;
        RECT 25.104 20.544 25.136 21.288 ;
  LAYER M1 ;
        RECT 25.184 20.544 25.216 21.288 ;
  LAYER M1 ;
        RECT 25.184 21.384 25.216 21.624 ;
  LAYER M1 ;
        RECT 25.184 21.888 25.216 22.128 ;
  LAYER M1 ;
        RECT 25.264 20.544 25.296 21.288 ;
  LAYER M1 ;
        RECT 25.344 20.544 25.376 21.288 ;
  LAYER M1 ;
        RECT 25.344 21.384 25.376 21.624 ;
  LAYER M1 ;
        RECT 25.344 21.888 25.376 22.128 ;
  LAYER M1 ;
        RECT 25.424 20.544 25.456 21.288 ;
  LAYER M1 ;
        RECT 25.504 20.544 25.536 21.288 ;
  LAYER M1 ;
        RECT 25.504 21.384 25.536 21.624 ;
  LAYER M1 ;
        RECT 25.504 21.888 25.536 22.128 ;
  LAYER M1 ;
        RECT 25.584 20.544 25.616 21.288 ;
  LAYER M1 ;
        RECT 25.664 20.544 25.696 21.288 ;
  LAYER M1 ;
        RECT 25.664 21.384 25.696 21.624 ;
  LAYER M1 ;
        RECT 25.664 21.888 25.696 22.128 ;
  LAYER M1 ;
        RECT 25.744 20.544 25.776 21.288 ;
  LAYER M1 ;
        RECT 25.824 20.544 25.856 21.288 ;
  LAYER M1 ;
        RECT 25.824 21.384 25.856 21.624 ;
  LAYER M1 ;
        RECT 25.824 21.888 25.856 22.128 ;
  LAYER M1 ;
        RECT 25.904 20.544 25.936 21.288 ;
  LAYER M1 ;
        RECT 25.984 20.544 26.016 21.288 ;
  LAYER M1 ;
        RECT 25.984 21.384 26.016 21.624 ;
  LAYER M1 ;
        RECT 25.984 21.888 26.016 22.128 ;
  LAYER M1 ;
        RECT 26.064 20.544 26.096 21.288 ;
  LAYER M1 ;
        RECT 26.144 20.544 26.176 21.288 ;
  LAYER M1 ;
        RECT 26.144 21.384 26.176 21.624 ;
  LAYER M1 ;
        RECT 26.144 21.888 26.176 22.128 ;
  LAYER M1 ;
        RECT 26.224 20.544 26.256 21.288 ;
  LAYER M1 ;
        RECT 26.304 20.544 26.336 21.288 ;
  LAYER M1 ;
        RECT 26.304 21.384 26.336 21.624 ;
  LAYER M1 ;
        RECT 26.304 21.888 26.336 22.128 ;
  LAYER M1 ;
        RECT 26.384 20.544 26.416 21.288 ;
  LAYER M1 ;
        RECT 26.464 20.544 26.496 21.288 ;
  LAYER M1 ;
        RECT 26.464 21.384 26.496 21.624 ;
  LAYER M1 ;
        RECT 26.464 21.888 26.496 22.128 ;
  LAYER M1 ;
        RECT 26.544 20.544 26.576 21.288 ;
  LAYER M1 ;
        RECT 26.624 20.544 26.656 21.288 ;
  LAYER M1 ;
        RECT 26.624 21.384 26.656 21.624 ;
  LAYER M1 ;
        RECT 26.624 21.888 26.656 22.128 ;
  LAYER M1 ;
        RECT 26.704 20.544 26.736 21.288 ;
  LAYER M1 ;
        RECT 26.784 20.544 26.816 21.288 ;
  LAYER M1 ;
        RECT 26.784 21.384 26.816 21.624 ;
  LAYER M1 ;
        RECT 26.784 21.888 26.816 22.128 ;
  LAYER M1 ;
        RECT 26.864 20.544 26.896 21.288 ;
  LAYER M1 ;
        RECT 26.944 20.544 26.976 21.288 ;
  LAYER M1 ;
        RECT 26.944 21.384 26.976 21.624 ;
  LAYER M1 ;
        RECT 26.944 21.888 26.976 22.128 ;
  LAYER M1 ;
        RECT 27.024 20.544 27.056 21.288 ;
  LAYER M1 ;
        RECT 7.344 18.612 7.376 19.356 ;
  LAYER M1 ;
        RECT 7.344 19.452 7.376 19.692 ;
  LAYER M1 ;
        RECT 7.344 19.956 7.376 20.196 ;
  LAYER M1 ;
        RECT 7.264 18.612 7.296 19.356 ;
  LAYER M1 ;
        RECT 7.424 18.612 7.456 19.356 ;
  LAYER M1 ;
        RECT 7.504 18.612 7.536 19.356 ;
  LAYER M1 ;
        RECT 7.504 19.452 7.536 19.692 ;
  LAYER M1 ;
        RECT 7.504 19.956 7.536 20.196 ;
  LAYER M1 ;
        RECT 7.584 18.612 7.616 19.356 ;
  LAYER M1 ;
        RECT 7.664 18.612 7.696 19.356 ;
  LAYER M1 ;
        RECT 7.664 19.452 7.696 19.692 ;
  LAYER M1 ;
        RECT 7.664 19.956 7.696 20.196 ;
  LAYER M1 ;
        RECT 7.744 18.612 7.776 19.356 ;
  LAYER M1 ;
        RECT 7.824 18.612 7.856 19.356 ;
  LAYER M1 ;
        RECT 7.824 19.452 7.856 19.692 ;
  LAYER M1 ;
        RECT 7.824 19.956 7.856 20.196 ;
  LAYER M1 ;
        RECT 7.904 18.612 7.936 19.356 ;
  LAYER M1 ;
        RECT 7.984 18.612 8.016 19.356 ;
  LAYER M1 ;
        RECT 7.984 19.452 8.016 19.692 ;
  LAYER M1 ;
        RECT 7.984 19.956 8.016 20.196 ;
  LAYER M1 ;
        RECT 8.064 18.612 8.096 19.356 ;
  LAYER M1 ;
        RECT 8.144 18.612 8.176 19.356 ;
  LAYER M1 ;
        RECT 8.144 19.452 8.176 19.692 ;
  LAYER M1 ;
        RECT 8.144 19.956 8.176 20.196 ;
  LAYER M1 ;
        RECT 8.224 18.612 8.256 19.356 ;
  LAYER M1 ;
        RECT 8.304 18.612 8.336 19.356 ;
  LAYER M1 ;
        RECT 8.304 19.452 8.336 19.692 ;
  LAYER M1 ;
        RECT 8.304 19.956 8.336 20.196 ;
  LAYER M1 ;
        RECT 8.384 18.612 8.416 19.356 ;
  LAYER M1 ;
        RECT 8.464 18.612 8.496 19.356 ;
  LAYER M1 ;
        RECT 8.464 19.452 8.496 19.692 ;
  LAYER M1 ;
        RECT 8.464 19.956 8.496 20.196 ;
  LAYER M1 ;
        RECT 8.544 18.612 8.576 19.356 ;
  LAYER M1 ;
        RECT 8.624 18.612 8.656 19.356 ;
  LAYER M1 ;
        RECT 8.624 19.452 8.656 19.692 ;
  LAYER M1 ;
        RECT 8.624 19.956 8.656 20.196 ;
  LAYER M1 ;
        RECT 8.704 18.612 8.736 19.356 ;
  LAYER M1 ;
        RECT 8.784 18.612 8.816 19.356 ;
  LAYER M1 ;
        RECT 8.784 19.452 8.816 19.692 ;
  LAYER M1 ;
        RECT 8.784 19.956 8.816 20.196 ;
  LAYER M1 ;
        RECT 8.864 18.612 8.896 19.356 ;
  LAYER M1 ;
        RECT 8.944 18.612 8.976 19.356 ;
  LAYER M1 ;
        RECT 8.944 19.452 8.976 19.692 ;
  LAYER M1 ;
        RECT 8.944 19.956 8.976 20.196 ;
  LAYER M1 ;
        RECT 9.024 18.612 9.056 19.356 ;
  LAYER M1 ;
        RECT 9.104 18.612 9.136 19.356 ;
  LAYER M1 ;
        RECT 9.104 19.452 9.136 19.692 ;
  LAYER M1 ;
        RECT 9.104 19.956 9.136 20.196 ;
  LAYER M1 ;
        RECT 9.184 18.612 9.216 19.356 ;
  LAYER M1 ;
        RECT 9.264 18.612 9.296 19.356 ;
  LAYER M1 ;
        RECT 9.264 19.452 9.296 19.692 ;
  LAYER M1 ;
        RECT 9.264 19.956 9.296 20.196 ;
  LAYER M1 ;
        RECT 9.344 18.612 9.376 19.356 ;
  LAYER M1 ;
        RECT 9.424 18.612 9.456 19.356 ;
  LAYER M1 ;
        RECT 9.424 19.452 9.456 19.692 ;
  LAYER M1 ;
        RECT 9.424 19.956 9.456 20.196 ;
  LAYER M1 ;
        RECT 9.504 18.612 9.536 19.356 ;
  LAYER M1 ;
        RECT 9.584 18.612 9.616 19.356 ;
  LAYER M1 ;
        RECT 9.584 19.452 9.616 19.692 ;
  LAYER M1 ;
        RECT 9.584 19.956 9.616 20.196 ;
  LAYER M1 ;
        RECT 9.664 18.612 9.696 19.356 ;
  LAYER M1 ;
        RECT 9.744 18.612 9.776 19.356 ;
  LAYER M1 ;
        RECT 9.744 19.452 9.776 19.692 ;
  LAYER M1 ;
        RECT 9.744 19.956 9.776 20.196 ;
  LAYER M1 ;
        RECT 9.824 18.612 9.856 19.356 ;
  LAYER M1 ;
        RECT 9.904 18.612 9.936 19.356 ;
  LAYER M1 ;
        RECT 9.904 19.452 9.936 19.692 ;
  LAYER M1 ;
        RECT 9.904 19.956 9.936 20.196 ;
  LAYER M1 ;
        RECT 9.984 18.612 10.016 19.356 ;
  LAYER M1 ;
        RECT 10.064 18.612 10.096 19.356 ;
  LAYER M1 ;
        RECT 10.064 19.452 10.096 19.692 ;
  LAYER M1 ;
        RECT 10.064 19.956 10.096 20.196 ;
  LAYER M1 ;
        RECT 10.144 18.612 10.176 19.356 ;
  LAYER M1 ;
        RECT 10.224 18.612 10.256 19.356 ;
  LAYER M1 ;
        RECT 10.224 19.452 10.256 19.692 ;
  LAYER M1 ;
        RECT 10.224 19.956 10.256 20.196 ;
  LAYER M1 ;
        RECT 10.304 18.612 10.336 19.356 ;
  LAYER M1 ;
        RECT 10.384 18.612 10.416 19.356 ;
  LAYER M1 ;
        RECT 10.384 19.452 10.416 19.692 ;
  LAYER M1 ;
        RECT 10.384 19.956 10.416 20.196 ;
  LAYER M1 ;
        RECT 10.464 18.612 10.496 19.356 ;
  LAYER M1 ;
        RECT 10.544 18.612 10.576 19.356 ;
  LAYER M1 ;
        RECT 10.544 19.452 10.576 19.692 ;
  LAYER M1 ;
        RECT 10.544 19.956 10.576 20.196 ;
  LAYER M1 ;
        RECT 10.624 18.612 10.656 19.356 ;
  LAYER M1 ;
        RECT 10.704 18.612 10.736 19.356 ;
  LAYER M1 ;
        RECT 10.704 19.452 10.736 19.692 ;
  LAYER M1 ;
        RECT 10.704 19.956 10.736 20.196 ;
  LAYER M1 ;
        RECT 10.784 18.612 10.816 19.356 ;
  LAYER M1 ;
        RECT 10.864 18.612 10.896 19.356 ;
  LAYER M1 ;
        RECT 10.864 19.452 10.896 19.692 ;
  LAYER M1 ;
        RECT 10.864 19.956 10.896 20.196 ;
  LAYER M1 ;
        RECT 10.944 18.612 10.976 19.356 ;
  LAYER M1 ;
        RECT 11.024 18.612 11.056 19.356 ;
  LAYER M1 ;
        RECT 11.024 19.452 11.056 19.692 ;
  LAYER M1 ;
        RECT 11.024 19.956 11.056 20.196 ;
  LAYER M1 ;
        RECT 11.104 18.612 11.136 19.356 ;
  LAYER M1 ;
        RECT 11.184 18.612 11.216 19.356 ;
  LAYER M1 ;
        RECT 11.184 19.452 11.216 19.692 ;
  LAYER M1 ;
        RECT 11.184 19.956 11.216 20.196 ;
  LAYER M1 ;
        RECT 11.264 18.612 11.296 19.356 ;
  LAYER M1 ;
        RECT 11.344 18.612 11.376 19.356 ;
  LAYER M1 ;
        RECT 11.344 19.452 11.376 19.692 ;
  LAYER M1 ;
        RECT 11.344 19.956 11.376 20.196 ;
  LAYER M1 ;
        RECT 11.424 18.612 11.456 19.356 ;
  LAYER M1 ;
        RECT 11.504 18.612 11.536 19.356 ;
  LAYER M1 ;
        RECT 11.504 19.452 11.536 19.692 ;
  LAYER M1 ;
        RECT 11.504 19.956 11.536 20.196 ;
  LAYER M1 ;
        RECT 11.584 18.612 11.616 19.356 ;
  LAYER M1 ;
        RECT 11.664 18.612 11.696 19.356 ;
  LAYER M1 ;
        RECT 11.664 19.452 11.696 19.692 ;
  LAYER M1 ;
        RECT 11.664 19.956 11.696 20.196 ;
  LAYER M1 ;
        RECT 11.744 18.612 11.776 19.356 ;
  LAYER M1 ;
        RECT 11.824 18.612 11.856 19.356 ;
  LAYER M1 ;
        RECT 11.824 19.452 11.856 19.692 ;
  LAYER M1 ;
        RECT 11.824 19.956 11.856 20.196 ;
  LAYER M1 ;
        RECT 11.904 18.612 11.936 19.356 ;
  LAYER M1 ;
        RECT 11.984 18.612 12.016 19.356 ;
  LAYER M1 ;
        RECT 11.984 19.452 12.016 19.692 ;
  LAYER M1 ;
        RECT 11.984 19.956 12.016 20.196 ;
  LAYER M1 ;
        RECT 12.064 18.612 12.096 19.356 ;
  LAYER M1 ;
        RECT 12.144 18.612 12.176 19.356 ;
  LAYER M1 ;
        RECT 12.144 19.452 12.176 19.692 ;
  LAYER M1 ;
        RECT 12.144 19.956 12.176 20.196 ;
  LAYER M1 ;
        RECT 12.224 18.612 12.256 19.356 ;
  LAYER M1 ;
        RECT 12.304 18.612 12.336 19.356 ;
  LAYER M1 ;
        RECT 12.304 19.452 12.336 19.692 ;
  LAYER M1 ;
        RECT 12.304 19.956 12.336 20.196 ;
  LAYER M1 ;
        RECT 12.384 18.612 12.416 19.356 ;
  LAYER M1 ;
        RECT 12.464 18.612 12.496 19.356 ;
  LAYER M1 ;
        RECT 12.464 19.452 12.496 19.692 ;
  LAYER M1 ;
        RECT 12.464 19.956 12.496 20.196 ;
  LAYER M1 ;
        RECT 12.544 18.612 12.576 19.356 ;
  LAYER M1 ;
        RECT 12.624 18.612 12.656 19.356 ;
  LAYER M1 ;
        RECT 12.624 19.452 12.656 19.692 ;
  LAYER M1 ;
        RECT 12.624 19.956 12.656 20.196 ;
  LAYER M1 ;
        RECT 12.704 18.612 12.736 19.356 ;
  LAYER M1 ;
        RECT 12.784 18.612 12.816 19.356 ;
  LAYER M1 ;
        RECT 12.784 19.452 12.816 19.692 ;
  LAYER M1 ;
        RECT 12.784 19.956 12.816 20.196 ;
  LAYER M1 ;
        RECT 12.864 18.612 12.896 19.356 ;
  LAYER M1 ;
        RECT 12.944 18.612 12.976 19.356 ;
  LAYER M1 ;
        RECT 12.944 19.452 12.976 19.692 ;
  LAYER M1 ;
        RECT 12.944 19.956 12.976 20.196 ;
  LAYER M1 ;
        RECT 13.024 18.612 13.056 19.356 ;
  LAYER M1 ;
        RECT 13.104 18.612 13.136 19.356 ;
  LAYER M1 ;
        RECT 13.104 19.452 13.136 19.692 ;
  LAYER M1 ;
        RECT 13.104 19.956 13.136 20.196 ;
  LAYER M1 ;
        RECT 13.184 18.612 13.216 19.356 ;
  LAYER M1 ;
        RECT 13.264 18.612 13.296 19.356 ;
  LAYER M1 ;
        RECT 13.264 19.452 13.296 19.692 ;
  LAYER M1 ;
        RECT 13.264 19.956 13.296 20.196 ;
  LAYER M1 ;
        RECT 13.344 18.612 13.376 19.356 ;
  LAYER M1 ;
        RECT 13.424 18.612 13.456 19.356 ;
  LAYER M1 ;
        RECT 13.424 19.452 13.456 19.692 ;
  LAYER M1 ;
        RECT 13.424 19.956 13.456 20.196 ;
  LAYER M1 ;
        RECT 13.504 18.612 13.536 19.356 ;
  LAYER M1 ;
        RECT 13.584 18.612 13.616 19.356 ;
  LAYER M1 ;
        RECT 13.584 19.452 13.616 19.692 ;
  LAYER M1 ;
        RECT 13.584 19.956 13.616 20.196 ;
  LAYER M1 ;
        RECT 13.664 18.612 13.696 19.356 ;
  LAYER M1 ;
        RECT 13.744 18.612 13.776 19.356 ;
  LAYER M1 ;
        RECT 13.744 19.452 13.776 19.692 ;
  LAYER M1 ;
        RECT 13.744 19.956 13.776 20.196 ;
  LAYER M1 ;
        RECT 13.824 18.612 13.856 19.356 ;
  LAYER M1 ;
        RECT 13.904 18.612 13.936 19.356 ;
  LAYER M1 ;
        RECT 13.904 19.452 13.936 19.692 ;
  LAYER M1 ;
        RECT 13.904 19.956 13.936 20.196 ;
  LAYER M1 ;
        RECT 13.984 18.612 14.016 19.356 ;
  LAYER M1 ;
        RECT 14.064 18.612 14.096 19.356 ;
  LAYER M1 ;
        RECT 14.064 19.452 14.096 19.692 ;
  LAYER M1 ;
        RECT 14.064 19.956 14.096 20.196 ;
  LAYER M1 ;
        RECT 14.144 18.612 14.176 19.356 ;
  LAYER M1 ;
        RECT 14.224 18.612 14.256 19.356 ;
  LAYER M1 ;
        RECT 14.224 19.452 14.256 19.692 ;
  LAYER M1 ;
        RECT 14.224 19.956 14.256 20.196 ;
  LAYER M1 ;
        RECT 14.304 18.612 14.336 19.356 ;
  LAYER M1 ;
        RECT 14.384 18.612 14.416 19.356 ;
  LAYER M1 ;
        RECT 14.384 19.452 14.416 19.692 ;
  LAYER M1 ;
        RECT 14.384 19.956 14.416 20.196 ;
  LAYER M1 ;
        RECT 14.464 18.612 14.496 19.356 ;
  LAYER M1 ;
        RECT 14.544 18.612 14.576 19.356 ;
  LAYER M1 ;
        RECT 14.544 19.452 14.576 19.692 ;
  LAYER M1 ;
        RECT 14.544 19.956 14.576 20.196 ;
  LAYER M1 ;
        RECT 14.624 18.612 14.656 19.356 ;
  LAYER M1 ;
        RECT 14.704 18.612 14.736 19.356 ;
  LAYER M1 ;
        RECT 14.704 19.452 14.736 19.692 ;
  LAYER M1 ;
        RECT 14.704 19.956 14.736 20.196 ;
  LAYER M1 ;
        RECT 14.784 18.612 14.816 19.356 ;
  LAYER M1 ;
        RECT 14.864 18.612 14.896 19.356 ;
  LAYER M1 ;
        RECT 14.864 19.452 14.896 19.692 ;
  LAYER M1 ;
        RECT 14.864 19.956 14.896 20.196 ;
  LAYER M1 ;
        RECT 14.944 18.612 14.976 19.356 ;
  LAYER M1 ;
        RECT 15.024 18.612 15.056 19.356 ;
  LAYER M1 ;
        RECT 15.024 19.452 15.056 19.692 ;
  LAYER M1 ;
        RECT 15.024 19.956 15.056 20.196 ;
  LAYER M1 ;
        RECT 15.104 18.612 15.136 19.356 ;
  LAYER M1 ;
        RECT 15.184 18.612 15.216 19.356 ;
  LAYER M1 ;
        RECT 15.184 19.452 15.216 19.692 ;
  LAYER M1 ;
        RECT 15.184 19.956 15.216 20.196 ;
  LAYER M1 ;
        RECT 15.264 18.612 15.296 19.356 ;
  LAYER M1 ;
        RECT 15.344 18.612 15.376 19.356 ;
  LAYER M1 ;
        RECT 15.344 19.452 15.376 19.692 ;
  LAYER M1 ;
        RECT 15.344 19.956 15.376 20.196 ;
  LAYER M1 ;
        RECT 15.424 18.612 15.456 19.356 ;
  LAYER M1 ;
        RECT 15.504 18.612 15.536 19.356 ;
  LAYER M1 ;
        RECT 15.504 19.452 15.536 19.692 ;
  LAYER M1 ;
        RECT 15.504 19.956 15.536 20.196 ;
  LAYER M1 ;
        RECT 15.584 18.612 15.616 19.356 ;
  LAYER M1 ;
        RECT 15.664 18.612 15.696 19.356 ;
  LAYER M1 ;
        RECT 15.664 19.452 15.696 19.692 ;
  LAYER M1 ;
        RECT 15.664 19.956 15.696 20.196 ;
  LAYER M1 ;
        RECT 15.744 18.612 15.776 19.356 ;
  LAYER M1 ;
        RECT 15.824 18.612 15.856 19.356 ;
  LAYER M1 ;
        RECT 15.824 19.452 15.856 19.692 ;
  LAYER M1 ;
        RECT 15.824 19.956 15.856 20.196 ;
  LAYER M1 ;
        RECT 15.904 18.612 15.936 19.356 ;
  LAYER M1 ;
        RECT 15.984 18.612 16.016 19.356 ;
  LAYER M1 ;
        RECT 15.984 19.452 16.016 19.692 ;
  LAYER M1 ;
        RECT 15.984 19.956 16.016 20.196 ;
  LAYER M1 ;
        RECT 16.064 18.612 16.096 19.356 ;
  LAYER M1 ;
        RECT 16.144 18.612 16.176 19.356 ;
  LAYER M1 ;
        RECT 16.144 19.452 16.176 19.692 ;
  LAYER M1 ;
        RECT 16.144 19.956 16.176 20.196 ;
  LAYER M1 ;
        RECT 16.224 18.612 16.256 19.356 ;
  LAYER M1 ;
        RECT 16.304 18.612 16.336 19.356 ;
  LAYER M1 ;
        RECT 16.304 19.452 16.336 19.692 ;
  LAYER M1 ;
        RECT 16.304 19.956 16.336 20.196 ;
  LAYER M1 ;
        RECT 16.384 18.612 16.416 19.356 ;
  LAYER M1 ;
        RECT 16.464 18.612 16.496 19.356 ;
  LAYER M1 ;
        RECT 16.464 19.452 16.496 19.692 ;
  LAYER M1 ;
        RECT 16.464 19.956 16.496 20.196 ;
  LAYER M1 ;
        RECT 16.544 18.612 16.576 19.356 ;
  LAYER M1 ;
        RECT 16.624 18.612 16.656 19.356 ;
  LAYER M1 ;
        RECT 16.624 19.452 16.656 19.692 ;
  LAYER M1 ;
        RECT 16.624 19.956 16.656 20.196 ;
  LAYER M1 ;
        RECT 16.704 18.612 16.736 19.356 ;
  LAYER M1 ;
        RECT 16.784 18.612 16.816 19.356 ;
  LAYER M1 ;
        RECT 16.784 19.452 16.816 19.692 ;
  LAYER M1 ;
        RECT 16.784 19.956 16.816 20.196 ;
  LAYER M1 ;
        RECT 16.864 18.612 16.896 19.356 ;
  LAYER M1 ;
        RECT 16.944 18.612 16.976 19.356 ;
  LAYER M1 ;
        RECT 16.944 19.452 16.976 19.692 ;
  LAYER M1 ;
        RECT 16.944 19.956 16.976 20.196 ;
  LAYER M1 ;
        RECT 17.024 18.612 17.056 19.356 ;
  LAYER M1 ;
        RECT 17.104 18.612 17.136 19.356 ;
  LAYER M1 ;
        RECT 17.104 19.452 17.136 19.692 ;
  LAYER M1 ;
        RECT 17.104 19.956 17.136 20.196 ;
  LAYER M1 ;
        RECT 17.184 18.612 17.216 19.356 ;
  LAYER M1 ;
        RECT 17.264 18.612 17.296 19.356 ;
  LAYER M1 ;
        RECT 17.264 19.452 17.296 19.692 ;
  LAYER M1 ;
        RECT 17.264 19.956 17.296 20.196 ;
  LAYER M1 ;
        RECT 17.344 18.612 17.376 19.356 ;
  LAYER M1 ;
        RECT 17.424 18.612 17.456 19.356 ;
  LAYER M1 ;
        RECT 17.424 19.452 17.456 19.692 ;
  LAYER M1 ;
        RECT 17.424 19.956 17.456 20.196 ;
  LAYER M1 ;
        RECT 17.504 18.612 17.536 19.356 ;
  LAYER M1 ;
        RECT 17.584 18.612 17.616 19.356 ;
  LAYER M1 ;
        RECT 17.584 19.452 17.616 19.692 ;
  LAYER M1 ;
        RECT 17.584 19.956 17.616 20.196 ;
  LAYER M1 ;
        RECT 17.664 18.612 17.696 19.356 ;
  LAYER M1 ;
        RECT 17.744 18.612 17.776 19.356 ;
  LAYER M1 ;
        RECT 17.744 19.452 17.776 19.692 ;
  LAYER M1 ;
        RECT 17.744 19.956 17.776 20.196 ;
  LAYER M1 ;
        RECT 17.824 18.612 17.856 19.356 ;
  LAYER M1 ;
        RECT 17.904 18.612 17.936 19.356 ;
  LAYER M1 ;
        RECT 17.904 19.452 17.936 19.692 ;
  LAYER M1 ;
        RECT 17.904 19.956 17.936 20.196 ;
  LAYER M1 ;
        RECT 17.984 18.612 18.016 19.356 ;
  LAYER M1 ;
        RECT 27.664 0.132 27.696 0.876 ;
  LAYER M1 ;
        RECT 27.664 0.972 27.696 1.212 ;
  LAYER M1 ;
        RECT 27.664 1.308 27.696 2.052 ;
  LAYER M1 ;
        RECT 27.664 2.148 27.696 2.388 ;
  LAYER M1 ;
        RECT 27.664 2.484 27.696 3.228 ;
  LAYER M1 ;
        RECT 27.664 3.324 27.696 3.564 ;
  LAYER M1 ;
        RECT 27.664 3.66 27.696 4.404 ;
  LAYER M1 ;
        RECT 27.664 4.5 27.696 4.74 ;
  LAYER M1 ;
        RECT 27.664 4.836 27.696 5.58 ;
  LAYER M1 ;
        RECT 27.664 5.676 27.696 5.916 ;
  LAYER M1 ;
        RECT 27.664 6.012 27.696 6.756 ;
  LAYER M1 ;
        RECT 27.664 6.852 27.696 7.092 ;
  LAYER M1 ;
        RECT 27.664 7.188 27.696 7.932 ;
  LAYER M1 ;
        RECT 27.664 8.028 27.696 8.268 ;
  LAYER M1 ;
        RECT 27.664 8.364 27.696 9.108 ;
  LAYER M1 ;
        RECT 27.664 9.204 27.696 9.444 ;
  LAYER M1 ;
        RECT 27.664 9.54 27.696 10.284 ;
  LAYER M1 ;
        RECT 27.664 10.38 27.696 10.62 ;
  LAYER M1 ;
        RECT 27.664 10.716 27.696 11.46 ;
  LAYER M1 ;
        RECT 27.664 11.556 27.696 11.796 ;
  LAYER M1 ;
        RECT 27.664 12.06 27.696 12.3 ;
  LAYER M1 ;
        RECT 27.584 0.132 27.616 0.876 ;
  LAYER M1 ;
        RECT 27.584 1.308 27.616 2.052 ;
  LAYER M1 ;
        RECT 27.584 2.484 27.616 3.228 ;
  LAYER M1 ;
        RECT 27.584 3.66 27.616 4.404 ;
  LAYER M1 ;
        RECT 27.584 4.836 27.616 5.58 ;
  LAYER M1 ;
        RECT 27.584 6.012 27.616 6.756 ;
  LAYER M1 ;
        RECT 27.584 7.188 27.616 7.932 ;
  LAYER M1 ;
        RECT 27.584 8.364 27.616 9.108 ;
  LAYER M1 ;
        RECT 27.584 9.54 27.616 10.284 ;
  LAYER M1 ;
        RECT 27.584 10.716 27.616 11.46 ;
  LAYER M1 ;
        RECT 27.744 0.132 27.776 0.876 ;
  LAYER M1 ;
        RECT 27.744 1.308 27.776 2.052 ;
  LAYER M1 ;
        RECT 27.744 2.484 27.776 3.228 ;
  LAYER M1 ;
        RECT 27.744 3.66 27.776 4.404 ;
  LAYER M1 ;
        RECT 27.744 4.836 27.776 5.58 ;
  LAYER M1 ;
        RECT 27.744 6.012 27.776 6.756 ;
  LAYER M1 ;
        RECT 27.744 7.188 27.776 7.932 ;
  LAYER M1 ;
        RECT 27.744 8.364 27.776 9.108 ;
  LAYER M1 ;
        RECT 27.744 9.54 27.776 10.284 ;
  LAYER M1 ;
        RECT 27.744 10.716 27.776 11.46 ;
  LAYER M1 ;
        RECT 27.824 0.132 27.856 0.876 ;
  LAYER M1 ;
        RECT 27.824 0.972 27.856 1.212 ;
  LAYER M1 ;
        RECT 27.824 1.308 27.856 2.052 ;
  LAYER M1 ;
        RECT 27.824 2.148 27.856 2.388 ;
  LAYER M1 ;
        RECT 27.824 2.484 27.856 3.228 ;
  LAYER M1 ;
        RECT 27.824 3.324 27.856 3.564 ;
  LAYER M1 ;
        RECT 27.824 3.66 27.856 4.404 ;
  LAYER M1 ;
        RECT 27.824 4.5 27.856 4.74 ;
  LAYER M1 ;
        RECT 27.824 4.836 27.856 5.58 ;
  LAYER M1 ;
        RECT 27.824 5.676 27.856 5.916 ;
  LAYER M1 ;
        RECT 27.824 6.012 27.856 6.756 ;
  LAYER M1 ;
        RECT 27.824 6.852 27.856 7.092 ;
  LAYER M1 ;
        RECT 27.824 7.188 27.856 7.932 ;
  LAYER M1 ;
        RECT 27.824 8.028 27.856 8.268 ;
  LAYER M1 ;
        RECT 27.824 8.364 27.856 9.108 ;
  LAYER M1 ;
        RECT 27.824 9.204 27.856 9.444 ;
  LAYER M1 ;
        RECT 27.824 9.54 27.856 10.284 ;
  LAYER M1 ;
        RECT 27.824 10.38 27.856 10.62 ;
  LAYER M1 ;
        RECT 27.824 10.716 27.856 11.46 ;
  LAYER M1 ;
        RECT 27.824 11.556 27.856 11.796 ;
  LAYER M1 ;
        RECT 27.824 12.06 27.856 12.3 ;
  LAYER M1 ;
        RECT 27.904 0.132 27.936 0.876 ;
  LAYER M1 ;
        RECT 27.904 1.308 27.936 2.052 ;
  LAYER M1 ;
        RECT 27.904 2.484 27.936 3.228 ;
  LAYER M1 ;
        RECT 27.904 3.66 27.936 4.404 ;
  LAYER M1 ;
        RECT 27.904 4.836 27.936 5.58 ;
  LAYER M1 ;
        RECT 27.904 6.012 27.936 6.756 ;
  LAYER M1 ;
        RECT 27.904 7.188 27.936 7.932 ;
  LAYER M1 ;
        RECT 27.904 8.364 27.936 9.108 ;
  LAYER M1 ;
        RECT 27.904 9.54 27.936 10.284 ;
  LAYER M1 ;
        RECT 27.904 10.716 27.936 11.46 ;
  LAYER M1 ;
        RECT 27.984 0.132 28.016 0.876 ;
  LAYER M1 ;
        RECT 27.984 0.972 28.016 1.212 ;
  LAYER M1 ;
        RECT 27.984 1.308 28.016 2.052 ;
  LAYER M1 ;
        RECT 27.984 2.148 28.016 2.388 ;
  LAYER M1 ;
        RECT 27.984 2.484 28.016 3.228 ;
  LAYER M1 ;
        RECT 27.984 3.324 28.016 3.564 ;
  LAYER M1 ;
        RECT 27.984 3.66 28.016 4.404 ;
  LAYER M1 ;
        RECT 27.984 4.5 28.016 4.74 ;
  LAYER M1 ;
        RECT 27.984 4.836 28.016 5.58 ;
  LAYER M1 ;
        RECT 27.984 5.676 28.016 5.916 ;
  LAYER M1 ;
        RECT 27.984 6.012 28.016 6.756 ;
  LAYER M1 ;
        RECT 27.984 6.852 28.016 7.092 ;
  LAYER M1 ;
        RECT 27.984 7.188 28.016 7.932 ;
  LAYER M1 ;
        RECT 27.984 8.028 28.016 8.268 ;
  LAYER M1 ;
        RECT 27.984 8.364 28.016 9.108 ;
  LAYER M1 ;
        RECT 27.984 9.204 28.016 9.444 ;
  LAYER M1 ;
        RECT 27.984 9.54 28.016 10.284 ;
  LAYER M1 ;
        RECT 27.984 10.38 28.016 10.62 ;
  LAYER M1 ;
        RECT 27.984 10.716 28.016 11.46 ;
  LAYER M1 ;
        RECT 27.984 11.556 28.016 11.796 ;
  LAYER M1 ;
        RECT 27.984 12.06 28.016 12.3 ;
  LAYER M1 ;
        RECT 28.064 0.132 28.096 0.876 ;
  LAYER M1 ;
        RECT 28.064 1.308 28.096 2.052 ;
  LAYER M1 ;
        RECT 28.064 2.484 28.096 3.228 ;
  LAYER M1 ;
        RECT 28.064 3.66 28.096 4.404 ;
  LAYER M1 ;
        RECT 28.064 4.836 28.096 5.58 ;
  LAYER M1 ;
        RECT 28.064 6.012 28.096 6.756 ;
  LAYER M1 ;
        RECT 28.064 7.188 28.096 7.932 ;
  LAYER M1 ;
        RECT 28.064 8.364 28.096 9.108 ;
  LAYER M1 ;
        RECT 28.064 9.54 28.096 10.284 ;
  LAYER M1 ;
        RECT 28.064 10.716 28.096 11.46 ;
  LAYER M1 ;
        RECT 28.144 0.132 28.176 0.876 ;
  LAYER M1 ;
        RECT 28.144 0.972 28.176 1.212 ;
  LAYER M1 ;
        RECT 28.144 1.308 28.176 2.052 ;
  LAYER M1 ;
        RECT 28.144 2.148 28.176 2.388 ;
  LAYER M1 ;
        RECT 28.144 2.484 28.176 3.228 ;
  LAYER M1 ;
        RECT 28.144 3.324 28.176 3.564 ;
  LAYER M1 ;
        RECT 28.144 3.66 28.176 4.404 ;
  LAYER M1 ;
        RECT 28.144 4.5 28.176 4.74 ;
  LAYER M1 ;
        RECT 28.144 4.836 28.176 5.58 ;
  LAYER M1 ;
        RECT 28.144 5.676 28.176 5.916 ;
  LAYER M1 ;
        RECT 28.144 6.012 28.176 6.756 ;
  LAYER M1 ;
        RECT 28.144 6.852 28.176 7.092 ;
  LAYER M1 ;
        RECT 28.144 7.188 28.176 7.932 ;
  LAYER M1 ;
        RECT 28.144 8.028 28.176 8.268 ;
  LAYER M1 ;
        RECT 28.144 8.364 28.176 9.108 ;
  LAYER M1 ;
        RECT 28.144 9.204 28.176 9.444 ;
  LAYER M1 ;
        RECT 28.144 9.54 28.176 10.284 ;
  LAYER M1 ;
        RECT 28.144 10.38 28.176 10.62 ;
  LAYER M1 ;
        RECT 28.144 10.716 28.176 11.46 ;
  LAYER M1 ;
        RECT 28.144 11.556 28.176 11.796 ;
  LAYER M1 ;
        RECT 28.144 12.06 28.176 12.3 ;
  LAYER M1 ;
        RECT 28.224 0.132 28.256 0.876 ;
  LAYER M1 ;
        RECT 28.224 1.308 28.256 2.052 ;
  LAYER M1 ;
        RECT 28.224 2.484 28.256 3.228 ;
  LAYER M1 ;
        RECT 28.224 3.66 28.256 4.404 ;
  LAYER M1 ;
        RECT 28.224 4.836 28.256 5.58 ;
  LAYER M1 ;
        RECT 28.224 6.012 28.256 6.756 ;
  LAYER M1 ;
        RECT 28.224 7.188 28.256 7.932 ;
  LAYER M1 ;
        RECT 28.224 8.364 28.256 9.108 ;
  LAYER M1 ;
        RECT 28.224 9.54 28.256 10.284 ;
  LAYER M1 ;
        RECT 28.224 10.716 28.256 11.46 ;
  LAYER M1 ;
        RECT 28.304 0.132 28.336 0.876 ;
  LAYER M1 ;
        RECT 28.304 0.972 28.336 1.212 ;
  LAYER M1 ;
        RECT 28.304 1.308 28.336 2.052 ;
  LAYER M1 ;
        RECT 28.304 2.148 28.336 2.388 ;
  LAYER M1 ;
        RECT 28.304 2.484 28.336 3.228 ;
  LAYER M1 ;
        RECT 28.304 3.324 28.336 3.564 ;
  LAYER M1 ;
        RECT 28.304 3.66 28.336 4.404 ;
  LAYER M1 ;
        RECT 28.304 4.5 28.336 4.74 ;
  LAYER M1 ;
        RECT 28.304 4.836 28.336 5.58 ;
  LAYER M1 ;
        RECT 28.304 5.676 28.336 5.916 ;
  LAYER M1 ;
        RECT 28.304 6.012 28.336 6.756 ;
  LAYER M1 ;
        RECT 28.304 6.852 28.336 7.092 ;
  LAYER M1 ;
        RECT 28.304 7.188 28.336 7.932 ;
  LAYER M1 ;
        RECT 28.304 8.028 28.336 8.268 ;
  LAYER M1 ;
        RECT 28.304 8.364 28.336 9.108 ;
  LAYER M1 ;
        RECT 28.304 9.204 28.336 9.444 ;
  LAYER M1 ;
        RECT 28.304 9.54 28.336 10.284 ;
  LAYER M1 ;
        RECT 28.304 10.38 28.336 10.62 ;
  LAYER M1 ;
        RECT 28.304 10.716 28.336 11.46 ;
  LAYER M1 ;
        RECT 28.304 11.556 28.336 11.796 ;
  LAYER M1 ;
        RECT 28.304 12.06 28.336 12.3 ;
  LAYER M1 ;
        RECT 28.384 0.132 28.416 0.876 ;
  LAYER M1 ;
        RECT 28.384 1.308 28.416 2.052 ;
  LAYER M1 ;
        RECT 28.384 2.484 28.416 3.228 ;
  LAYER M1 ;
        RECT 28.384 3.66 28.416 4.404 ;
  LAYER M1 ;
        RECT 28.384 4.836 28.416 5.58 ;
  LAYER M1 ;
        RECT 28.384 6.012 28.416 6.756 ;
  LAYER M1 ;
        RECT 28.384 7.188 28.416 7.932 ;
  LAYER M1 ;
        RECT 28.384 8.364 28.416 9.108 ;
  LAYER M1 ;
        RECT 28.384 9.54 28.416 10.284 ;
  LAYER M1 ;
        RECT 28.384 10.716 28.416 11.46 ;
  LAYER M1 ;
        RECT 28.464 0.132 28.496 0.876 ;
  LAYER M1 ;
        RECT 28.464 0.972 28.496 1.212 ;
  LAYER M1 ;
        RECT 28.464 1.308 28.496 2.052 ;
  LAYER M1 ;
        RECT 28.464 2.148 28.496 2.388 ;
  LAYER M1 ;
        RECT 28.464 2.484 28.496 3.228 ;
  LAYER M1 ;
        RECT 28.464 3.324 28.496 3.564 ;
  LAYER M1 ;
        RECT 28.464 3.66 28.496 4.404 ;
  LAYER M1 ;
        RECT 28.464 4.5 28.496 4.74 ;
  LAYER M1 ;
        RECT 28.464 4.836 28.496 5.58 ;
  LAYER M1 ;
        RECT 28.464 5.676 28.496 5.916 ;
  LAYER M1 ;
        RECT 28.464 6.012 28.496 6.756 ;
  LAYER M1 ;
        RECT 28.464 6.852 28.496 7.092 ;
  LAYER M1 ;
        RECT 28.464 7.188 28.496 7.932 ;
  LAYER M1 ;
        RECT 28.464 8.028 28.496 8.268 ;
  LAYER M1 ;
        RECT 28.464 8.364 28.496 9.108 ;
  LAYER M1 ;
        RECT 28.464 9.204 28.496 9.444 ;
  LAYER M1 ;
        RECT 28.464 9.54 28.496 10.284 ;
  LAYER M1 ;
        RECT 28.464 10.38 28.496 10.62 ;
  LAYER M1 ;
        RECT 28.464 10.716 28.496 11.46 ;
  LAYER M1 ;
        RECT 28.464 11.556 28.496 11.796 ;
  LAYER M1 ;
        RECT 28.464 12.06 28.496 12.3 ;
  LAYER M1 ;
        RECT 28.544 0.132 28.576 0.876 ;
  LAYER M1 ;
        RECT 28.544 1.308 28.576 2.052 ;
  LAYER M1 ;
        RECT 28.544 2.484 28.576 3.228 ;
  LAYER M1 ;
        RECT 28.544 3.66 28.576 4.404 ;
  LAYER M1 ;
        RECT 28.544 4.836 28.576 5.58 ;
  LAYER M1 ;
        RECT 28.544 6.012 28.576 6.756 ;
  LAYER M1 ;
        RECT 28.544 7.188 28.576 7.932 ;
  LAYER M1 ;
        RECT 28.544 8.364 28.576 9.108 ;
  LAYER M1 ;
        RECT 28.544 9.54 28.576 10.284 ;
  LAYER M1 ;
        RECT 28.544 10.716 28.576 11.46 ;
  LAYER M1 ;
        RECT 28.624 0.132 28.656 0.876 ;
  LAYER M1 ;
        RECT 28.624 0.972 28.656 1.212 ;
  LAYER M1 ;
        RECT 28.624 1.308 28.656 2.052 ;
  LAYER M1 ;
        RECT 28.624 2.148 28.656 2.388 ;
  LAYER M1 ;
        RECT 28.624 2.484 28.656 3.228 ;
  LAYER M1 ;
        RECT 28.624 3.324 28.656 3.564 ;
  LAYER M1 ;
        RECT 28.624 3.66 28.656 4.404 ;
  LAYER M1 ;
        RECT 28.624 4.5 28.656 4.74 ;
  LAYER M1 ;
        RECT 28.624 4.836 28.656 5.58 ;
  LAYER M1 ;
        RECT 28.624 5.676 28.656 5.916 ;
  LAYER M1 ;
        RECT 28.624 6.012 28.656 6.756 ;
  LAYER M1 ;
        RECT 28.624 6.852 28.656 7.092 ;
  LAYER M1 ;
        RECT 28.624 7.188 28.656 7.932 ;
  LAYER M1 ;
        RECT 28.624 8.028 28.656 8.268 ;
  LAYER M1 ;
        RECT 28.624 8.364 28.656 9.108 ;
  LAYER M1 ;
        RECT 28.624 9.204 28.656 9.444 ;
  LAYER M1 ;
        RECT 28.624 9.54 28.656 10.284 ;
  LAYER M1 ;
        RECT 28.624 10.38 28.656 10.62 ;
  LAYER M1 ;
        RECT 28.624 10.716 28.656 11.46 ;
  LAYER M1 ;
        RECT 28.624 11.556 28.656 11.796 ;
  LAYER M1 ;
        RECT 28.624 12.06 28.656 12.3 ;
  LAYER M1 ;
        RECT 28.704 0.132 28.736 0.876 ;
  LAYER M1 ;
        RECT 28.704 1.308 28.736 2.052 ;
  LAYER M1 ;
        RECT 28.704 2.484 28.736 3.228 ;
  LAYER M1 ;
        RECT 28.704 3.66 28.736 4.404 ;
  LAYER M1 ;
        RECT 28.704 4.836 28.736 5.58 ;
  LAYER M1 ;
        RECT 28.704 6.012 28.736 6.756 ;
  LAYER M1 ;
        RECT 28.704 7.188 28.736 7.932 ;
  LAYER M1 ;
        RECT 28.704 8.364 28.736 9.108 ;
  LAYER M1 ;
        RECT 28.704 9.54 28.736 10.284 ;
  LAYER M1 ;
        RECT 28.704 10.716 28.736 11.46 ;
  LAYER M1 ;
        RECT 28.784 0.132 28.816 0.876 ;
  LAYER M1 ;
        RECT 28.784 0.972 28.816 1.212 ;
  LAYER M1 ;
        RECT 28.784 1.308 28.816 2.052 ;
  LAYER M1 ;
        RECT 28.784 2.148 28.816 2.388 ;
  LAYER M1 ;
        RECT 28.784 2.484 28.816 3.228 ;
  LAYER M1 ;
        RECT 28.784 3.324 28.816 3.564 ;
  LAYER M1 ;
        RECT 28.784 3.66 28.816 4.404 ;
  LAYER M1 ;
        RECT 28.784 4.5 28.816 4.74 ;
  LAYER M1 ;
        RECT 28.784 4.836 28.816 5.58 ;
  LAYER M1 ;
        RECT 28.784 5.676 28.816 5.916 ;
  LAYER M1 ;
        RECT 28.784 6.012 28.816 6.756 ;
  LAYER M1 ;
        RECT 28.784 6.852 28.816 7.092 ;
  LAYER M1 ;
        RECT 28.784 7.188 28.816 7.932 ;
  LAYER M1 ;
        RECT 28.784 8.028 28.816 8.268 ;
  LAYER M1 ;
        RECT 28.784 8.364 28.816 9.108 ;
  LAYER M1 ;
        RECT 28.784 9.204 28.816 9.444 ;
  LAYER M1 ;
        RECT 28.784 9.54 28.816 10.284 ;
  LAYER M1 ;
        RECT 28.784 10.38 28.816 10.62 ;
  LAYER M1 ;
        RECT 28.784 10.716 28.816 11.46 ;
  LAYER M1 ;
        RECT 28.784 11.556 28.816 11.796 ;
  LAYER M1 ;
        RECT 28.784 12.06 28.816 12.3 ;
  LAYER M1 ;
        RECT 28.864 0.132 28.896 0.876 ;
  LAYER M1 ;
        RECT 28.864 1.308 28.896 2.052 ;
  LAYER M1 ;
        RECT 28.864 2.484 28.896 3.228 ;
  LAYER M1 ;
        RECT 28.864 3.66 28.896 4.404 ;
  LAYER M1 ;
        RECT 28.864 4.836 28.896 5.58 ;
  LAYER M1 ;
        RECT 28.864 6.012 28.896 6.756 ;
  LAYER M1 ;
        RECT 28.864 7.188 28.896 7.932 ;
  LAYER M1 ;
        RECT 28.864 8.364 28.896 9.108 ;
  LAYER M1 ;
        RECT 28.864 9.54 28.896 10.284 ;
  LAYER M1 ;
        RECT 28.864 10.716 28.896 11.46 ;
  LAYER M1 ;
        RECT 28.944 0.132 28.976 0.876 ;
  LAYER M1 ;
        RECT 28.944 0.972 28.976 1.212 ;
  LAYER M1 ;
        RECT 28.944 1.308 28.976 2.052 ;
  LAYER M1 ;
        RECT 28.944 2.148 28.976 2.388 ;
  LAYER M1 ;
        RECT 28.944 2.484 28.976 3.228 ;
  LAYER M1 ;
        RECT 28.944 3.324 28.976 3.564 ;
  LAYER M1 ;
        RECT 28.944 3.66 28.976 4.404 ;
  LAYER M1 ;
        RECT 28.944 4.5 28.976 4.74 ;
  LAYER M1 ;
        RECT 28.944 4.836 28.976 5.58 ;
  LAYER M1 ;
        RECT 28.944 5.676 28.976 5.916 ;
  LAYER M1 ;
        RECT 28.944 6.012 28.976 6.756 ;
  LAYER M1 ;
        RECT 28.944 6.852 28.976 7.092 ;
  LAYER M1 ;
        RECT 28.944 7.188 28.976 7.932 ;
  LAYER M1 ;
        RECT 28.944 8.028 28.976 8.268 ;
  LAYER M1 ;
        RECT 28.944 8.364 28.976 9.108 ;
  LAYER M1 ;
        RECT 28.944 9.204 28.976 9.444 ;
  LAYER M1 ;
        RECT 28.944 9.54 28.976 10.284 ;
  LAYER M1 ;
        RECT 28.944 10.38 28.976 10.62 ;
  LAYER M1 ;
        RECT 28.944 10.716 28.976 11.46 ;
  LAYER M1 ;
        RECT 28.944 11.556 28.976 11.796 ;
  LAYER M1 ;
        RECT 28.944 12.06 28.976 12.3 ;
  LAYER M1 ;
        RECT 29.024 0.132 29.056 0.876 ;
  LAYER M1 ;
        RECT 29.024 1.308 29.056 2.052 ;
  LAYER M1 ;
        RECT 29.024 2.484 29.056 3.228 ;
  LAYER M1 ;
        RECT 29.024 3.66 29.056 4.404 ;
  LAYER M1 ;
        RECT 29.024 4.836 29.056 5.58 ;
  LAYER M1 ;
        RECT 29.024 6.012 29.056 6.756 ;
  LAYER M1 ;
        RECT 29.024 7.188 29.056 7.932 ;
  LAYER M1 ;
        RECT 29.024 8.364 29.056 9.108 ;
  LAYER M1 ;
        RECT 29.024 9.54 29.056 10.284 ;
  LAYER M1 ;
        RECT 29.024 10.716 29.056 11.46 ;
  LAYER M1 ;
        RECT 29.104 0.132 29.136 0.876 ;
  LAYER M1 ;
        RECT 29.104 0.972 29.136 1.212 ;
  LAYER M1 ;
        RECT 29.104 1.308 29.136 2.052 ;
  LAYER M1 ;
        RECT 29.104 2.148 29.136 2.388 ;
  LAYER M1 ;
        RECT 29.104 2.484 29.136 3.228 ;
  LAYER M1 ;
        RECT 29.104 3.324 29.136 3.564 ;
  LAYER M1 ;
        RECT 29.104 3.66 29.136 4.404 ;
  LAYER M1 ;
        RECT 29.104 4.5 29.136 4.74 ;
  LAYER M1 ;
        RECT 29.104 4.836 29.136 5.58 ;
  LAYER M1 ;
        RECT 29.104 5.676 29.136 5.916 ;
  LAYER M1 ;
        RECT 29.104 6.012 29.136 6.756 ;
  LAYER M1 ;
        RECT 29.104 6.852 29.136 7.092 ;
  LAYER M1 ;
        RECT 29.104 7.188 29.136 7.932 ;
  LAYER M1 ;
        RECT 29.104 8.028 29.136 8.268 ;
  LAYER M1 ;
        RECT 29.104 8.364 29.136 9.108 ;
  LAYER M1 ;
        RECT 29.104 9.204 29.136 9.444 ;
  LAYER M1 ;
        RECT 29.104 9.54 29.136 10.284 ;
  LAYER M1 ;
        RECT 29.104 10.38 29.136 10.62 ;
  LAYER M1 ;
        RECT 29.104 10.716 29.136 11.46 ;
  LAYER M1 ;
        RECT 29.104 11.556 29.136 11.796 ;
  LAYER M1 ;
        RECT 29.104 12.06 29.136 12.3 ;
  LAYER M1 ;
        RECT 29.184 0.132 29.216 0.876 ;
  LAYER M1 ;
        RECT 29.184 1.308 29.216 2.052 ;
  LAYER M1 ;
        RECT 29.184 2.484 29.216 3.228 ;
  LAYER M1 ;
        RECT 29.184 3.66 29.216 4.404 ;
  LAYER M1 ;
        RECT 29.184 4.836 29.216 5.58 ;
  LAYER M1 ;
        RECT 29.184 6.012 29.216 6.756 ;
  LAYER M1 ;
        RECT 29.184 7.188 29.216 7.932 ;
  LAYER M1 ;
        RECT 29.184 8.364 29.216 9.108 ;
  LAYER M1 ;
        RECT 29.184 9.54 29.216 10.284 ;
  LAYER M1 ;
        RECT 29.184 10.716 29.216 11.46 ;
  LAYER M1 ;
        RECT 29.264 0.132 29.296 0.876 ;
  LAYER M1 ;
        RECT 29.264 0.972 29.296 1.212 ;
  LAYER M1 ;
        RECT 29.264 1.308 29.296 2.052 ;
  LAYER M1 ;
        RECT 29.264 2.148 29.296 2.388 ;
  LAYER M1 ;
        RECT 29.264 2.484 29.296 3.228 ;
  LAYER M1 ;
        RECT 29.264 3.324 29.296 3.564 ;
  LAYER M1 ;
        RECT 29.264 3.66 29.296 4.404 ;
  LAYER M1 ;
        RECT 29.264 4.5 29.296 4.74 ;
  LAYER M1 ;
        RECT 29.264 4.836 29.296 5.58 ;
  LAYER M1 ;
        RECT 29.264 5.676 29.296 5.916 ;
  LAYER M1 ;
        RECT 29.264 6.012 29.296 6.756 ;
  LAYER M1 ;
        RECT 29.264 6.852 29.296 7.092 ;
  LAYER M1 ;
        RECT 29.264 7.188 29.296 7.932 ;
  LAYER M1 ;
        RECT 29.264 8.028 29.296 8.268 ;
  LAYER M1 ;
        RECT 29.264 8.364 29.296 9.108 ;
  LAYER M1 ;
        RECT 29.264 9.204 29.296 9.444 ;
  LAYER M1 ;
        RECT 29.264 9.54 29.296 10.284 ;
  LAYER M1 ;
        RECT 29.264 10.38 29.296 10.62 ;
  LAYER M1 ;
        RECT 29.264 10.716 29.296 11.46 ;
  LAYER M1 ;
        RECT 29.264 11.556 29.296 11.796 ;
  LAYER M1 ;
        RECT 29.264 12.06 29.296 12.3 ;
  LAYER M1 ;
        RECT 29.344 0.132 29.376 0.876 ;
  LAYER M1 ;
        RECT 29.344 1.308 29.376 2.052 ;
  LAYER M1 ;
        RECT 29.344 2.484 29.376 3.228 ;
  LAYER M1 ;
        RECT 29.344 3.66 29.376 4.404 ;
  LAYER M1 ;
        RECT 29.344 4.836 29.376 5.58 ;
  LAYER M1 ;
        RECT 29.344 6.012 29.376 6.756 ;
  LAYER M1 ;
        RECT 29.344 7.188 29.376 7.932 ;
  LAYER M1 ;
        RECT 29.344 8.364 29.376 9.108 ;
  LAYER M1 ;
        RECT 29.344 9.54 29.376 10.284 ;
  LAYER M1 ;
        RECT 29.344 10.716 29.376 11.46 ;
  LAYER M1 ;
        RECT 29.424 0.132 29.456 0.876 ;
  LAYER M1 ;
        RECT 29.424 0.972 29.456 1.212 ;
  LAYER M1 ;
        RECT 29.424 1.308 29.456 2.052 ;
  LAYER M1 ;
        RECT 29.424 2.148 29.456 2.388 ;
  LAYER M1 ;
        RECT 29.424 2.484 29.456 3.228 ;
  LAYER M1 ;
        RECT 29.424 3.324 29.456 3.564 ;
  LAYER M1 ;
        RECT 29.424 3.66 29.456 4.404 ;
  LAYER M1 ;
        RECT 29.424 4.5 29.456 4.74 ;
  LAYER M1 ;
        RECT 29.424 4.836 29.456 5.58 ;
  LAYER M1 ;
        RECT 29.424 5.676 29.456 5.916 ;
  LAYER M1 ;
        RECT 29.424 6.012 29.456 6.756 ;
  LAYER M1 ;
        RECT 29.424 6.852 29.456 7.092 ;
  LAYER M1 ;
        RECT 29.424 7.188 29.456 7.932 ;
  LAYER M1 ;
        RECT 29.424 8.028 29.456 8.268 ;
  LAYER M1 ;
        RECT 29.424 8.364 29.456 9.108 ;
  LAYER M1 ;
        RECT 29.424 9.204 29.456 9.444 ;
  LAYER M1 ;
        RECT 29.424 9.54 29.456 10.284 ;
  LAYER M1 ;
        RECT 29.424 10.38 29.456 10.62 ;
  LAYER M1 ;
        RECT 29.424 10.716 29.456 11.46 ;
  LAYER M1 ;
        RECT 29.424 11.556 29.456 11.796 ;
  LAYER M1 ;
        RECT 29.424 12.06 29.456 12.3 ;
  LAYER M1 ;
        RECT 29.504 0.132 29.536 0.876 ;
  LAYER M1 ;
        RECT 29.504 1.308 29.536 2.052 ;
  LAYER M1 ;
        RECT 29.504 2.484 29.536 3.228 ;
  LAYER M1 ;
        RECT 29.504 3.66 29.536 4.404 ;
  LAYER M1 ;
        RECT 29.504 4.836 29.536 5.58 ;
  LAYER M1 ;
        RECT 29.504 6.012 29.536 6.756 ;
  LAYER M1 ;
        RECT 29.504 7.188 29.536 7.932 ;
  LAYER M1 ;
        RECT 29.504 8.364 29.536 9.108 ;
  LAYER M1 ;
        RECT 29.504 9.54 29.536 10.284 ;
  LAYER M1 ;
        RECT 29.504 10.716 29.536 11.46 ;
  LAYER M1 ;
        RECT 29.584 0.132 29.616 0.876 ;
  LAYER M1 ;
        RECT 29.584 0.972 29.616 1.212 ;
  LAYER M1 ;
        RECT 29.584 1.308 29.616 2.052 ;
  LAYER M1 ;
        RECT 29.584 2.148 29.616 2.388 ;
  LAYER M1 ;
        RECT 29.584 2.484 29.616 3.228 ;
  LAYER M1 ;
        RECT 29.584 3.324 29.616 3.564 ;
  LAYER M1 ;
        RECT 29.584 3.66 29.616 4.404 ;
  LAYER M1 ;
        RECT 29.584 4.5 29.616 4.74 ;
  LAYER M1 ;
        RECT 29.584 4.836 29.616 5.58 ;
  LAYER M1 ;
        RECT 29.584 5.676 29.616 5.916 ;
  LAYER M1 ;
        RECT 29.584 6.012 29.616 6.756 ;
  LAYER M1 ;
        RECT 29.584 6.852 29.616 7.092 ;
  LAYER M1 ;
        RECT 29.584 7.188 29.616 7.932 ;
  LAYER M1 ;
        RECT 29.584 8.028 29.616 8.268 ;
  LAYER M1 ;
        RECT 29.584 8.364 29.616 9.108 ;
  LAYER M1 ;
        RECT 29.584 9.204 29.616 9.444 ;
  LAYER M1 ;
        RECT 29.584 9.54 29.616 10.284 ;
  LAYER M1 ;
        RECT 29.584 10.38 29.616 10.62 ;
  LAYER M1 ;
        RECT 29.584 10.716 29.616 11.46 ;
  LAYER M1 ;
        RECT 29.584 11.556 29.616 11.796 ;
  LAYER M1 ;
        RECT 29.584 12.06 29.616 12.3 ;
  LAYER M1 ;
        RECT 29.664 0.132 29.696 0.876 ;
  LAYER M1 ;
        RECT 29.664 1.308 29.696 2.052 ;
  LAYER M1 ;
        RECT 29.664 2.484 29.696 3.228 ;
  LAYER M1 ;
        RECT 29.664 3.66 29.696 4.404 ;
  LAYER M1 ;
        RECT 29.664 4.836 29.696 5.58 ;
  LAYER M1 ;
        RECT 29.664 6.012 29.696 6.756 ;
  LAYER M1 ;
        RECT 29.664 7.188 29.696 7.932 ;
  LAYER M1 ;
        RECT 29.664 8.364 29.696 9.108 ;
  LAYER M1 ;
        RECT 29.664 9.54 29.696 10.284 ;
  LAYER M1 ;
        RECT 29.664 10.716 29.696 11.46 ;
  LAYER M1 ;
        RECT 29.744 0.132 29.776 0.876 ;
  LAYER M1 ;
        RECT 29.744 0.972 29.776 1.212 ;
  LAYER M1 ;
        RECT 29.744 1.308 29.776 2.052 ;
  LAYER M1 ;
        RECT 29.744 2.148 29.776 2.388 ;
  LAYER M1 ;
        RECT 29.744 2.484 29.776 3.228 ;
  LAYER M1 ;
        RECT 29.744 3.324 29.776 3.564 ;
  LAYER M1 ;
        RECT 29.744 3.66 29.776 4.404 ;
  LAYER M1 ;
        RECT 29.744 4.5 29.776 4.74 ;
  LAYER M1 ;
        RECT 29.744 4.836 29.776 5.58 ;
  LAYER M1 ;
        RECT 29.744 5.676 29.776 5.916 ;
  LAYER M1 ;
        RECT 29.744 6.012 29.776 6.756 ;
  LAYER M1 ;
        RECT 29.744 6.852 29.776 7.092 ;
  LAYER M1 ;
        RECT 29.744 7.188 29.776 7.932 ;
  LAYER M1 ;
        RECT 29.744 8.028 29.776 8.268 ;
  LAYER M1 ;
        RECT 29.744 8.364 29.776 9.108 ;
  LAYER M1 ;
        RECT 29.744 9.204 29.776 9.444 ;
  LAYER M1 ;
        RECT 29.744 9.54 29.776 10.284 ;
  LAYER M1 ;
        RECT 29.744 10.38 29.776 10.62 ;
  LAYER M1 ;
        RECT 29.744 10.716 29.776 11.46 ;
  LAYER M1 ;
        RECT 29.744 11.556 29.776 11.796 ;
  LAYER M1 ;
        RECT 29.744 12.06 29.776 12.3 ;
  LAYER M1 ;
        RECT 29.824 0.132 29.856 0.876 ;
  LAYER M1 ;
        RECT 29.824 1.308 29.856 2.052 ;
  LAYER M1 ;
        RECT 29.824 2.484 29.856 3.228 ;
  LAYER M1 ;
        RECT 29.824 3.66 29.856 4.404 ;
  LAYER M1 ;
        RECT 29.824 4.836 29.856 5.58 ;
  LAYER M1 ;
        RECT 29.824 6.012 29.856 6.756 ;
  LAYER M1 ;
        RECT 29.824 7.188 29.856 7.932 ;
  LAYER M1 ;
        RECT 29.824 8.364 29.856 9.108 ;
  LAYER M1 ;
        RECT 29.824 9.54 29.856 10.284 ;
  LAYER M1 ;
        RECT 29.824 10.716 29.856 11.46 ;
  LAYER M1 ;
        RECT 29.904 0.132 29.936 0.876 ;
  LAYER M1 ;
        RECT 29.904 0.972 29.936 1.212 ;
  LAYER M1 ;
        RECT 29.904 1.308 29.936 2.052 ;
  LAYER M1 ;
        RECT 29.904 2.148 29.936 2.388 ;
  LAYER M1 ;
        RECT 29.904 2.484 29.936 3.228 ;
  LAYER M1 ;
        RECT 29.904 3.324 29.936 3.564 ;
  LAYER M1 ;
        RECT 29.904 3.66 29.936 4.404 ;
  LAYER M1 ;
        RECT 29.904 4.5 29.936 4.74 ;
  LAYER M1 ;
        RECT 29.904 4.836 29.936 5.58 ;
  LAYER M1 ;
        RECT 29.904 5.676 29.936 5.916 ;
  LAYER M1 ;
        RECT 29.904 6.012 29.936 6.756 ;
  LAYER M1 ;
        RECT 29.904 6.852 29.936 7.092 ;
  LAYER M1 ;
        RECT 29.904 7.188 29.936 7.932 ;
  LAYER M1 ;
        RECT 29.904 8.028 29.936 8.268 ;
  LAYER M1 ;
        RECT 29.904 8.364 29.936 9.108 ;
  LAYER M1 ;
        RECT 29.904 9.204 29.936 9.444 ;
  LAYER M1 ;
        RECT 29.904 9.54 29.936 10.284 ;
  LAYER M1 ;
        RECT 29.904 10.38 29.936 10.62 ;
  LAYER M1 ;
        RECT 29.904 10.716 29.936 11.46 ;
  LAYER M1 ;
        RECT 29.904 11.556 29.936 11.796 ;
  LAYER M1 ;
        RECT 29.904 12.06 29.936 12.3 ;
  LAYER M1 ;
        RECT 29.984 0.132 30.016 0.876 ;
  LAYER M1 ;
        RECT 29.984 1.308 30.016 2.052 ;
  LAYER M1 ;
        RECT 29.984 2.484 30.016 3.228 ;
  LAYER M1 ;
        RECT 29.984 3.66 30.016 4.404 ;
  LAYER M1 ;
        RECT 29.984 4.836 30.016 5.58 ;
  LAYER M1 ;
        RECT 29.984 6.012 30.016 6.756 ;
  LAYER M1 ;
        RECT 29.984 7.188 30.016 7.932 ;
  LAYER M1 ;
        RECT 29.984 8.364 30.016 9.108 ;
  LAYER M1 ;
        RECT 29.984 9.54 30.016 10.284 ;
  LAYER M1 ;
        RECT 29.984 10.716 30.016 11.46 ;
  LAYER M1 ;
        RECT 30.064 0.132 30.096 0.876 ;
  LAYER M1 ;
        RECT 30.064 0.972 30.096 1.212 ;
  LAYER M1 ;
        RECT 30.064 1.308 30.096 2.052 ;
  LAYER M1 ;
        RECT 30.064 2.148 30.096 2.388 ;
  LAYER M1 ;
        RECT 30.064 2.484 30.096 3.228 ;
  LAYER M1 ;
        RECT 30.064 3.324 30.096 3.564 ;
  LAYER M1 ;
        RECT 30.064 3.66 30.096 4.404 ;
  LAYER M1 ;
        RECT 30.064 4.5 30.096 4.74 ;
  LAYER M1 ;
        RECT 30.064 4.836 30.096 5.58 ;
  LAYER M1 ;
        RECT 30.064 5.676 30.096 5.916 ;
  LAYER M1 ;
        RECT 30.064 6.012 30.096 6.756 ;
  LAYER M1 ;
        RECT 30.064 6.852 30.096 7.092 ;
  LAYER M1 ;
        RECT 30.064 7.188 30.096 7.932 ;
  LAYER M1 ;
        RECT 30.064 8.028 30.096 8.268 ;
  LAYER M1 ;
        RECT 30.064 8.364 30.096 9.108 ;
  LAYER M1 ;
        RECT 30.064 9.204 30.096 9.444 ;
  LAYER M1 ;
        RECT 30.064 9.54 30.096 10.284 ;
  LAYER M1 ;
        RECT 30.064 10.38 30.096 10.62 ;
  LAYER M1 ;
        RECT 30.064 10.716 30.096 11.46 ;
  LAYER M1 ;
        RECT 30.064 11.556 30.096 11.796 ;
  LAYER M1 ;
        RECT 30.064 12.06 30.096 12.3 ;
  LAYER M1 ;
        RECT 30.144 0.132 30.176 0.876 ;
  LAYER M1 ;
        RECT 30.144 1.308 30.176 2.052 ;
  LAYER M1 ;
        RECT 30.144 2.484 30.176 3.228 ;
  LAYER M1 ;
        RECT 30.144 3.66 30.176 4.404 ;
  LAYER M1 ;
        RECT 30.144 4.836 30.176 5.58 ;
  LAYER M1 ;
        RECT 30.144 6.012 30.176 6.756 ;
  LAYER M1 ;
        RECT 30.144 7.188 30.176 7.932 ;
  LAYER M1 ;
        RECT 30.144 8.364 30.176 9.108 ;
  LAYER M1 ;
        RECT 30.144 9.54 30.176 10.284 ;
  LAYER M1 ;
        RECT 30.144 10.716 30.176 11.46 ;
  LAYER M1 ;
        RECT 30.224 0.132 30.256 0.876 ;
  LAYER M1 ;
        RECT 30.224 0.972 30.256 1.212 ;
  LAYER M1 ;
        RECT 30.224 1.308 30.256 2.052 ;
  LAYER M1 ;
        RECT 30.224 2.148 30.256 2.388 ;
  LAYER M1 ;
        RECT 30.224 2.484 30.256 3.228 ;
  LAYER M1 ;
        RECT 30.224 3.324 30.256 3.564 ;
  LAYER M1 ;
        RECT 30.224 3.66 30.256 4.404 ;
  LAYER M1 ;
        RECT 30.224 4.5 30.256 4.74 ;
  LAYER M1 ;
        RECT 30.224 4.836 30.256 5.58 ;
  LAYER M1 ;
        RECT 30.224 5.676 30.256 5.916 ;
  LAYER M1 ;
        RECT 30.224 6.012 30.256 6.756 ;
  LAYER M1 ;
        RECT 30.224 6.852 30.256 7.092 ;
  LAYER M1 ;
        RECT 30.224 7.188 30.256 7.932 ;
  LAYER M1 ;
        RECT 30.224 8.028 30.256 8.268 ;
  LAYER M1 ;
        RECT 30.224 8.364 30.256 9.108 ;
  LAYER M1 ;
        RECT 30.224 9.204 30.256 9.444 ;
  LAYER M1 ;
        RECT 30.224 9.54 30.256 10.284 ;
  LAYER M1 ;
        RECT 30.224 10.38 30.256 10.62 ;
  LAYER M1 ;
        RECT 30.224 10.716 30.256 11.46 ;
  LAYER M1 ;
        RECT 30.224 11.556 30.256 11.796 ;
  LAYER M1 ;
        RECT 30.224 12.06 30.256 12.3 ;
  LAYER M1 ;
        RECT 30.304 0.132 30.336 0.876 ;
  LAYER M1 ;
        RECT 30.304 1.308 30.336 2.052 ;
  LAYER M1 ;
        RECT 30.304 2.484 30.336 3.228 ;
  LAYER M1 ;
        RECT 30.304 3.66 30.336 4.404 ;
  LAYER M1 ;
        RECT 30.304 4.836 30.336 5.58 ;
  LAYER M1 ;
        RECT 30.304 6.012 30.336 6.756 ;
  LAYER M1 ;
        RECT 30.304 7.188 30.336 7.932 ;
  LAYER M1 ;
        RECT 30.304 8.364 30.336 9.108 ;
  LAYER M1 ;
        RECT 30.304 9.54 30.336 10.284 ;
  LAYER M1 ;
        RECT 30.304 10.716 30.336 11.46 ;
  LAYER M1 ;
        RECT 30.384 0.132 30.416 0.876 ;
  LAYER M1 ;
        RECT 30.384 0.972 30.416 1.212 ;
  LAYER M1 ;
        RECT 30.384 1.308 30.416 2.052 ;
  LAYER M1 ;
        RECT 30.384 2.148 30.416 2.388 ;
  LAYER M1 ;
        RECT 30.384 2.484 30.416 3.228 ;
  LAYER M1 ;
        RECT 30.384 3.324 30.416 3.564 ;
  LAYER M1 ;
        RECT 30.384 3.66 30.416 4.404 ;
  LAYER M1 ;
        RECT 30.384 4.5 30.416 4.74 ;
  LAYER M1 ;
        RECT 30.384 4.836 30.416 5.58 ;
  LAYER M1 ;
        RECT 30.384 5.676 30.416 5.916 ;
  LAYER M1 ;
        RECT 30.384 6.012 30.416 6.756 ;
  LAYER M1 ;
        RECT 30.384 6.852 30.416 7.092 ;
  LAYER M1 ;
        RECT 30.384 7.188 30.416 7.932 ;
  LAYER M1 ;
        RECT 30.384 8.028 30.416 8.268 ;
  LAYER M1 ;
        RECT 30.384 8.364 30.416 9.108 ;
  LAYER M1 ;
        RECT 30.384 9.204 30.416 9.444 ;
  LAYER M1 ;
        RECT 30.384 9.54 30.416 10.284 ;
  LAYER M1 ;
        RECT 30.384 10.38 30.416 10.62 ;
  LAYER M1 ;
        RECT 30.384 10.716 30.416 11.46 ;
  LAYER M1 ;
        RECT 30.384 11.556 30.416 11.796 ;
  LAYER M1 ;
        RECT 30.384 12.06 30.416 12.3 ;
  LAYER M1 ;
        RECT 30.464 0.132 30.496 0.876 ;
  LAYER M1 ;
        RECT 30.464 1.308 30.496 2.052 ;
  LAYER M1 ;
        RECT 30.464 2.484 30.496 3.228 ;
  LAYER M1 ;
        RECT 30.464 3.66 30.496 4.404 ;
  LAYER M1 ;
        RECT 30.464 4.836 30.496 5.58 ;
  LAYER M1 ;
        RECT 30.464 6.012 30.496 6.756 ;
  LAYER M1 ;
        RECT 30.464 7.188 30.496 7.932 ;
  LAYER M1 ;
        RECT 30.464 8.364 30.496 9.108 ;
  LAYER M1 ;
        RECT 30.464 9.54 30.496 10.284 ;
  LAYER M1 ;
        RECT 30.464 10.716 30.496 11.46 ;
  LAYER M1 ;
        RECT 30.544 0.132 30.576 0.876 ;
  LAYER M1 ;
        RECT 30.544 0.972 30.576 1.212 ;
  LAYER M1 ;
        RECT 30.544 1.308 30.576 2.052 ;
  LAYER M1 ;
        RECT 30.544 2.148 30.576 2.388 ;
  LAYER M1 ;
        RECT 30.544 2.484 30.576 3.228 ;
  LAYER M1 ;
        RECT 30.544 3.324 30.576 3.564 ;
  LAYER M1 ;
        RECT 30.544 3.66 30.576 4.404 ;
  LAYER M1 ;
        RECT 30.544 4.5 30.576 4.74 ;
  LAYER M1 ;
        RECT 30.544 4.836 30.576 5.58 ;
  LAYER M1 ;
        RECT 30.544 5.676 30.576 5.916 ;
  LAYER M1 ;
        RECT 30.544 6.012 30.576 6.756 ;
  LAYER M1 ;
        RECT 30.544 6.852 30.576 7.092 ;
  LAYER M1 ;
        RECT 30.544 7.188 30.576 7.932 ;
  LAYER M1 ;
        RECT 30.544 8.028 30.576 8.268 ;
  LAYER M1 ;
        RECT 30.544 8.364 30.576 9.108 ;
  LAYER M1 ;
        RECT 30.544 9.204 30.576 9.444 ;
  LAYER M1 ;
        RECT 30.544 9.54 30.576 10.284 ;
  LAYER M1 ;
        RECT 30.544 10.38 30.576 10.62 ;
  LAYER M1 ;
        RECT 30.544 10.716 30.576 11.46 ;
  LAYER M1 ;
        RECT 30.544 11.556 30.576 11.796 ;
  LAYER M1 ;
        RECT 30.544 12.06 30.576 12.3 ;
  LAYER M1 ;
        RECT 30.624 0.132 30.656 0.876 ;
  LAYER M1 ;
        RECT 30.624 1.308 30.656 2.052 ;
  LAYER M1 ;
        RECT 30.624 2.484 30.656 3.228 ;
  LAYER M1 ;
        RECT 30.624 3.66 30.656 4.404 ;
  LAYER M1 ;
        RECT 30.624 4.836 30.656 5.58 ;
  LAYER M1 ;
        RECT 30.624 6.012 30.656 6.756 ;
  LAYER M1 ;
        RECT 30.624 7.188 30.656 7.932 ;
  LAYER M1 ;
        RECT 30.624 8.364 30.656 9.108 ;
  LAYER M1 ;
        RECT 30.624 9.54 30.656 10.284 ;
  LAYER M1 ;
        RECT 30.624 10.716 30.656 11.46 ;
  LAYER M1 ;
        RECT 30.704 0.132 30.736 0.876 ;
  LAYER M1 ;
        RECT 30.704 0.972 30.736 1.212 ;
  LAYER M1 ;
        RECT 30.704 1.308 30.736 2.052 ;
  LAYER M1 ;
        RECT 30.704 2.148 30.736 2.388 ;
  LAYER M1 ;
        RECT 30.704 2.484 30.736 3.228 ;
  LAYER M1 ;
        RECT 30.704 3.324 30.736 3.564 ;
  LAYER M1 ;
        RECT 30.704 3.66 30.736 4.404 ;
  LAYER M1 ;
        RECT 30.704 4.5 30.736 4.74 ;
  LAYER M1 ;
        RECT 30.704 4.836 30.736 5.58 ;
  LAYER M1 ;
        RECT 30.704 5.676 30.736 5.916 ;
  LAYER M1 ;
        RECT 30.704 6.012 30.736 6.756 ;
  LAYER M1 ;
        RECT 30.704 6.852 30.736 7.092 ;
  LAYER M1 ;
        RECT 30.704 7.188 30.736 7.932 ;
  LAYER M1 ;
        RECT 30.704 8.028 30.736 8.268 ;
  LAYER M1 ;
        RECT 30.704 8.364 30.736 9.108 ;
  LAYER M1 ;
        RECT 30.704 9.204 30.736 9.444 ;
  LAYER M1 ;
        RECT 30.704 9.54 30.736 10.284 ;
  LAYER M1 ;
        RECT 30.704 10.38 30.736 10.62 ;
  LAYER M1 ;
        RECT 30.704 10.716 30.736 11.46 ;
  LAYER M1 ;
        RECT 30.704 11.556 30.736 11.796 ;
  LAYER M1 ;
        RECT 30.704 12.06 30.736 12.3 ;
  LAYER M1 ;
        RECT 30.784 0.132 30.816 0.876 ;
  LAYER M1 ;
        RECT 30.784 1.308 30.816 2.052 ;
  LAYER M1 ;
        RECT 30.784 2.484 30.816 3.228 ;
  LAYER M1 ;
        RECT 30.784 3.66 30.816 4.404 ;
  LAYER M1 ;
        RECT 30.784 4.836 30.816 5.58 ;
  LAYER M1 ;
        RECT 30.784 6.012 30.816 6.756 ;
  LAYER M1 ;
        RECT 30.784 7.188 30.816 7.932 ;
  LAYER M1 ;
        RECT 30.784 8.364 30.816 9.108 ;
  LAYER M1 ;
        RECT 30.784 9.54 30.816 10.284 ;
  LAYER M1 ;
        RECT 30.784 10.716 30.816 11.46 ;
  LAYER M1 ;
        RECT 30.864 0.132 30.896 0.876 ;
  LAYER M1 ;
        RECT 30.864 0.972 30.896 1.212 ;
  LAYER M1 ;
        RECT 30.864 1.308 30.896 2.052 ;
  LAYER M1 ;
        RECT 30.864 2.148 30.896 2.388 ;
  LAYER M1 ;
        RECT 30.864 2.484 30.896 3.228 ;
  LAYER M1 ;
        RECT 30.864 3.324 30.896 3.564 ;
  LAYER M1 ;
        RECT 30.864 3.66 30.896 4.404 ;
  LAYER M1 ;
        RECT 30.864 4.5 30.896 4.74 ;
  LAYER M1 ;
        RECT 30.864 4.836 30.896 5.58 ;
  LAYER M1 ;
        RECT 30.864 5.676 30.896 5.916 ;
  LAYER M1 ;
        RECT 30.864 6.012 30.896 6.756 ;
  LAYER M1 ;
        RECT 30.864 6.852 30.896 7.092 ;
  LAYER M1 ;
        RECT 30.864 7.188 30.896 7.932 ;
  LAYER M1 ;
        RECT 30.864 8.028 30.896 8.268 ;
  LAYER M1 ;
        RECT 30.864 8.364 30.896 9.108 ;
  LAYER M1 ;
        RECT 30.864 9.204 30.896 9.444 ;
  LAYER M1 ;
        RECT 30.864 9.54 30.896 10.284 ;
  LAYER M1 ;
        RECT 30.864 10.38 30.896 10.62 ;
  LAYER M1 ;
        RECT 30.864 10.716 30.896 11.46 ;
  LAYER M1 ;
        RECT 30.864 11.556 30.896 11.796 ;
  LAYER M1 ;
        RECT 30.864 12.06 30.896 12.3 ;
  LAYER M1 ;
        RECT 30.944 0.132 30.976 0.876 ;
  LAYER M1 ;
        RECT 30.944 1.308 30.976 2.052 ;
  LAYER M1 ;
        RECT 30.944 2.484 30.976 3.228 ;
  LAYER M1 ;
        RECT 30.944 3.66 30.976 4.404 ;
  LAYER M1 ;
        RECT 30.944 4.836 30.976 5.58 ;
  LAYER M1 ;
        RECT 30.944 6.012 30.976 6.756 ;
  LAYER M1 ;
        RECT 30.944 7.188 30.976 7.932 ;
  LAYER M1 ;
        RECT 30.944 8.364 30.976 9.108 ;
  LAYER M1 ;
        RECT 30.944 9.54 30.976 10.284 ;
  LAYER M1 ;
        RECT 30.944 10.716 30.976 11.46 ;
  LAYER M1 ;
        RECT 31.024 0.132 31.056 0.876 ;
  LAYER M1 ;
        RECT 31.024 0.972 31.056 1.212 ;
  LAYER M1 ;
        RECT 31.024 1.308 31.056 2.052 ;
  LAYER M1 ;
        RECT 31.024 2.148 31.056 2.388 ;
  LAYER M1 ;
        RECT 31.024 2.484 31.056 3.228 ;
  LAYER M1 ;
        RECT 31.024 3.324 31.056 3.564 ;
  LAYER M1 ;
        RECT 31.024 3.66 31.056 4.404 ;
  LAYER M1 ;
        RECT 31.024 4.5 31.056 4.74 ;
  LAYER M1 ;
        RECT 31.024 4.836 31.056 5.58 ;
  LAYER M1 ;
        RECT 31.024 5.676 31.056 5.916 ;
  LAYER M1 ;
        RECT 31.024 6.012 31.056 6.756 ;
  LAYER M1 ;
        RECT 31.024 6.852 31.056 7.092 ;
  LAYER M1 ;
        RECT 31.024 7.188 31.056 7.932 ;
  LAYER M1 ;
        RECT 31.024 8.028 31.056 8.268 ;
  LAYER M1 ;
        RECT 31.024 8.364 31.056 9.108 ;
  LAYER M1 ;
        RECT 31.024 9.204 31.056 9.444 ;
  LAYER M1 ;
        RECT 31.024 9.54 31.056 10.284 ;
  LAYER M1 ;
        RECT 31.024 10.38 31.056 10.62 ;
  LAYER M1 ;
        RECT 31.024 10.716 31.056 11.46 ;
  LAYER M1 ;
        RECT 31.024 11.556 31.056 11.796 ;
  LAYER M1 ;
        RECT 31.024 12.06 31.056 12.3 ;
  LAYER M1 ;
        RECT 31.104 0.132 31.136 0.876 ;
  LAYER M1 ;
        RECT 31.104 1.308 31.136 2.052 ;
  LAYER M1 ;
        RECT 31.104 2.484 31.136 3.228 ;
  LAYER M1 ;
        RECT 31.104 3.66 31.136 4.404 ;
  LAYER M1 ;
        RECT 31.104 4.836 31.136 5.58 ;
  LAYER M1 ;
        RECT 31.104 6.012 31.136 6.756 ;
  LAYER M1 ;
        RECT 31.104 7.188 31.136 7.932 ;
  LAYER M1 ;
        RECT 31.104 8.364 31.136 9.108 ;
  LAYER M1 ;
        RECT 31.104 9.54 31.136 10.284 ;
  LAYER M1 ;
        RECT 31.104 10.716 31.136 11.46 ;
  LAYER M1 ;
        RECT 31.184 0.132 31.216 0.876 ;
  LAYER M1 ;
        RECT 31.184 0.972 31.216 1.212 ;
  LAYER M1 ;
        RECT 31.184 1.308 31.216 2.052 ;
  LAYER M1 ;
        RECT 31.184 2.148 31.216 2.388 ;
  LAYER M1 ;
        RECT 31.184 2.484 31.216 3.228 ;
  LAYER M1 ;
        RECT 31.184 3.324 31.216 3.564 ;
  LAYER M1 ;
        RECT 31.184 3.66 31.216 4.404 ;
  LAYER M1 ;
        RECT 31.184 4.5 31.216 4.74 ;
  LAYER M1 ;
        RECT 31.184 4.836 31.216 5.58 ;
  LAYER M1 ;
        RECT 31.184 5.676 31.216 5.916 ;
  LAYER M1 ;
        RECT 31.184 6.012 31.216 6.756 ;
  LAYER M1 ;
        RECT 31.184 6.852 31.216 7.092 ;
  LAYER M1 ;
        RECT 31.184 7.188 31.216 7.932 ;
  LAYER M1 ;
        RECT 31.184 8.028 31.216 8.268 ;
  LAYER M1 ;
        RECT 31.184 8.364 31.216 9.108 ;
  LAYER M1 ;
        RECT 31.184 9.204 31.216 9.444 ;
  LAYER M1 ;
        RECT 31.184 9.54 31.216 10.284 ;
  LAYER M1 ;
        RECT 31.184 10.38 31.216 10.62 ;
  LAYER M1 ;
        RECT 31.184 10.716 31.216 11.46 ;
  LAYER M1 ;
        RECT 31.184 11.556 31.216 11.796 ;
  LAYER M1 ;
        RECT 31.184 12.06 31.216 12.3 ;
  LAYER M1 ;
        RECT 31.264 0.132 31.296 0.876 ;
  LAYER M1 ;
        RECT 31.264 1.308 31.296 2.052 ;
  LAYER M1 ;
        RECT 31.264 2.484 31.296 3.228 ;
  LAYER M1 ;
        RECT 31.264 3.66 31.296 4.404 ;
  LAYER M1 ;
        RECT 31.264 4.836 31.296 5.58 ;
  LAYER M1 ;
        RECT 31.264 6.012 31.296 6.756 ;
  LAYER M1 ;
        RECT 31.264 7.188 31.296 7.932 ;
  LAYER M1 ;
        RECT 31.264 8.364 31.296 9.108 ;
  LAYER M1 ;
        RECT 31.264 9.54 31.296 10.284 ;
  LAYER M1 ;
        RECT 31.264 10.716 31.296 11.46 ;
  LAYER M1 ;
        RECT 31.344 0.132 31.376 0.876 ;
  LAYER M1 ;
        RECT 31.344 0.972 31.376 1.212 ;
  LAYER M1 ;
        RECT 31.344 1.308 31.376 2.052 ;
  LAYER M1 ;
        RECT 31.344 2.148 31.376 2.388 ;
  LAYER M1 ;
        RECT 31.344 2.484 31.376 3.228 ;
  LAYER M1 ;
        RECT 31.344 3.324 31.376 3.564 ;
  LAYER M1 ;
        RECT 31.344 3.66 31.376 4.404 ;
  LAYER M1 ;
        RECT 31.344 4.5 31.376 4.74 ;
  LAYER M1 ;
        RECT 31.344 4.836 31.376 5.58 ;
  LAYER M1 ;
        RECT 31.344 5.676 31.376 5.916 ;
  LAYER M1 ;
        RECT 31.344 6.012 31.376 6.756 ;
  LAYER M1 ;
        RECT 31.344 6.852 31.376 7.092 ;
  LAYER M1 ;
        RECT 31.344 7.188 31.376 7.932 ;
  LAYER M1 ;
        RECT 31.344 8.028 31.376 8.268 ;
  LAYER M1 ;
        RECT 31.344 8.364 31.376 9.108 ;
  LAYER M1 ;
        RECT 31.344 9.204 31.376 9.444 ;
  LAYER M1 ;
        RECT 31.344 9.54 31.376 10.284 ;
  LAYER M1 ;
        RECT 31.344 10.38 31.376 10.62 ;
  LAYER M1 ;
        RECT 31.344 10.716 31.376 11.46 ;
  LAYER M1 ;
        RECT 31.344 11.556 31.376 11.796 ;
  LAYER M1 ;
        RECT 31.344 12.06 31.376 12.3 ;
  LAYER M1 ;
        RECT 31.424 0.132 31.456 0.876 ;
  LAYER M1 ;
        RECT 31.424 1.308 31.456 2.052 ;
  LAYER M1 ;
        RECT 31.424 2.484 31.456 3.228 ;
  LAYER M1 ;
        RECT 31.424 3.66 31.456 4.404 ;
  LAYER M1 ;
        RECT 31.424 4.836 31.456 5.58 ;
  LAYER M1 ;
        RECT 31.424 6.012 31.456 6.756 ;
  LAYER M1 ;
        RECT 31.424 7.188 31.456 7.932 ;
  LAYER M1 ;
        RECT 31.424 8.364 31.456 9.108 ;
  LAYER M1 ;
        RECT 31.424 9.54 31.456 10.284 ;
  LAYER M1 ;
        RECT 31.424 10.716 31.456 11.46 ;
  LAYER M1 ;
        RECT 31.504 0.132 31.536 0.876 ;
  LAYER M1 ;
        RECT 31.504 0.972 31.536 1.212 ;
  LAYER M1 ;
        RECT 31.504 1.308 31.536 2.052 ;
  LAYER M1 ;
        RECT 31.504 2.148 31.536 2.388 ;
  LAYER M1 ;
        RECT 31.504 2.484 31.536 3.228 ;
  LAYER M1 ;
        RECT 31.504 3.324 31.536 3.564 ;
  LAYER M1 ;
        RECT 31.504 3.66 31.536 4.404 ;
  LAYER M1 ;
        RECT 31.504 4.5 31.536 4.74 ;
  LAYER M1 ;
        RECT 31.504 4.836 31.536 5.58 ;
  LAYER M1 ;
        RECT 31.504 5.676 31.536 5.916 ;
  LAYER M1 ;
        RECT 31.504 6.012 31.536 6.756 ;
  LAYER M1 ;
        RECT 31.504 6.852 31.536 7.092 ;
  LAYER M1 ;
        RECT 31.504 7.188 31.536 7.932 ;
  LAYER M1 ;
        RECT 31.504 8.028 31.536 8.268 ;
  LAYER M1 ;
        RECT 31.504 8.364 31.536 9.108 ;
  LAYER M1 ;
        RECT 31.504 9.204 31.536 9.444 ;
  LAYER M1 ;
        RECT 31.504 9.54 31.536 10.284 ;
  LAYER M1 ;
        RECT 31.504 10.38 31.536 10.62 ;
  LAYER M1 ;
        RECT 31.504 10.716 31.536 11.46 ;
  LAYER M1 ;
        RECT 31.504 11.556 31.536 11.796 ;
  LAYER M1 ;
        RECT 31.504 12.06 31.536 12.3 ;
  LAYER M1 ;
        RECT 31.584 0.132 31.616 0.876 ;
  LAYER M1 ;
        RECT 31.584 1.308 31.616 2.052 ;
  LAYER M1 ;
        RECT 31.584 2.484 31.616 3.228 ;
  LAYER M1 ;
        RECT 31.584 3.66 31.616 4.404 ;
  LAYER M1 ;
        RECT 31.584 4.836 31.616 5.58 ;
  LAYER M1 ;
        RECT 31.584 6.012 31.616 6.756 ;
  LAYER M1 ;
        RECT 31.584 7.188 31.616 7.932 ;
  LAYER M1 ;
        RECT 31.584 8.364 31.616 9.108 ;
  LAYER M1 ;
        RECT 31.584 9.54 31.616 10.284 ;
  LAYER M1 ;
        RECT 31.584 10.716 31.616 11.46 ;
  LAYER M2 ;
        RECT 27.564 0.152 31.636 0.184 ;
  LAYER M2 ;
        RECT 27.644 0.236 31.556 0.268 ;
  LAYER M2 ;
        RECT 27.644 0.992 31.556 1.024 ;
  LAYER M2 ;
        RECT 27.564 1.328 31.636 1.36 ;
  LAYER M2 ;
        RECT 27.644 1.412 31.556 1.444 ;
  LAYER M2 ;
        RECT 27.644 2.168 31.556 2.2 ;
  LAYER M2 ;
        RECT 27.564 2.504 31.636 2.536 ;
  LAYER M2 ;
        RECT 27.644 2.588 31.556 2.62 ;
  LAYER M2 ;
        RECT 27.644 3.344 31.556 3.376 ;
  LAYER M2 ;
        RECT 27.564 3.68 31.636 3.712 ;
  LAYER M2 ;
        RECT 27.644 3.764 31.556 3.796 ;
  LAYER M2 ;
        RECT 27.644 4.52 31.556 4.552 ;
  LAYER M2 ;
        RECT 27.564 4.856 31.636 4.888 ;
  LAYER M2 ;
        RECT 27.644 4.94 31.556 4.972 ;
  LAYER M2 ;
        RECT 27.644 5.696 31.556 5.728 ;
  LAYER M2 ;
        RECT 27.564 6.032 31.636 6.064 ;
  LAYER M2 ;
        RECT 27.644 6.116 31.556 6.148 ;
  LAYER M2 ;
        RECT 27.644 6.872 31.556 6.904 ;
  LAYER M2 ;
        RECT 27.564 7.208 31.636 7.24 ;
  LAYER M2 ;
        RECT 27.644 7.292 31.556 7.324 ;
  LAYER M2 ;
        RECT 27.644 8.048 31.556 8.08 ;
  LAYER M2 ;
        RECT 27.564 8.384 31.636 8.416 ;
  LAYER M2 ;
        RECT 27.644 8.468 31.556 8.5 ;
  LAYER M2 ;
        RECT 27.644 9.224 31.556 9.256 ;
  LAYER M2 ;
        RECT 27.564 9.56 31.636 9.592 ;
  LAYER M2 ;
        RECT 27.644 9.644 31.556 9.676 ;
  LAYER M2 ;
        RECT 27.644 10.4 31.556 10.432 ;
  LAYER M2 ;
        RECT 27.564 10.736 31.636 10.768 ;
  LAYER M2 ;
        RECT 27.644 10.82 31.556 10.852 ;
  LAYER M2 ;
        RECT 27.644 11.576 31.556 11.608 ;
  LAYER M1 ;
        RECT 27.664 12.648 27.696 13.392 ;
  LAYER M1 ;
        RECT 27.664 13.488 27.696 13.728 ;
  LAYER M1 ;
        RECT 27.664 13.824 27.696 14.568 ;
  LAYER M1 ;
        RECT 27.664 14.664 27.696 14.904 ;
  LAYER M1 ;
        RECT 27.664 15 27.696 15.744 ;
  LAYER M1 ;
        RECT 27.664 15.84 27.696 16.08 ;
  LAYER M1 ;
        RECT 27.664 16.176 27.696 16.92 ;
  LAYER M1 ;
        RECT 27.664 17.016 27.696 17.256 ;
  LAYER M1 ;
        RECT 27.664 17.352 27.696 18.096 ;
  LAYER M1 ;
        RECT 27.664 18.192 27.696 18.432 ;
  LAYER M1 ;
        RECT 27.664 18.528 27.696 19.272 ;
  LAYER M1 ;
        RECT 27.664 19.368 27.696 19.608 ;
  LAYER M1 ;
        RECT 27.664 19.704 27.696 20.448 ;
  LAYER M1 ;
        RECT 27.664 20.544 27.696 20.784 ;
  LAYER M1 ;
        RECT 27.664 20.88 27.696 21.624 ;
  LAYER M1 ;
        RECT 27.664 21.72 27.696 21.96 ;
  LAYER M1 ;
        RECT 27.664 22.056 27.696 22.8 ;
  LAYER M1 ;
        RECT 27.664 22.896 27.696 23.136 ;
  LAYER M1 ;
        RECT 27.664 23.232 27.696 23.976 ;
  LAYER M1 ;
        RECT 27.664 24.072 27.696 24.312 ;
  LAYER M1 ;
        RECT 27.664 24.576 27.696 24.816 ;
  LAYER M1 ;
        RECT 27.584 12.648 27.616 13.392 ;
  LAYER M1 ;
        RECT 27.584 13.824 27.616 14.568 ;
  LAYER M1 ;
        RECT 27.584 15 27.616 15.744 ;
  LAYER M1 ;
        RECT 27.584 16.176 27.616 16.92 ;
  LAYER M1 ;
        RECT 27.584 17.352 27.616 18.096 ;
  LAYER M1 ;
        RECT 27.584 18.528 27.616 19.272 ;
  LAYER M1 ;
        RECT 27.584 19.704 27.616 20.448 ;
  LAYER M1 ;
        RECT 27.584 20.88 27.616 21.624 ;
  LAYER M1 ;
        RECT 27.584 22.056 27.616 22.8 ;
  LAYER M1 ;
        RECT 27.584 23.232 27.616 23.976 ;
  LAYER M1 ;
        RECT 27.744 12.648 27.776 13.392 ;
  LAYER M1 ;
        RECT 27.744 13.824 27.776 14.568 ;
  LAYER M1 ;
        RECT 27.744 15 27.776 15.744 ;
  LAYER M1 ;
        RECT 27.744 16.176 27.776 16.92 ;
  LAYER M1 ;
        RECT 27.744 17.352 27.776 18.096 ;
  LAYER M1 ;
        RECT 27.744 18.528 27.776 19.272 ;
  LAYER M1 ;
        RECT 27.744 19.704 27.776 20.448 ;
  LAYER M1 ;
        RECT 27.744 20.88 27.776 21.624 ;
  LAYER M1 ;
        RECT 27.744 22.056 27.776 22.8 ;
  LAYER M1 ;
        RECT 27.744 23.232 27.776 23.976 ;
  LAYER M1 ;
        RECT 27.824 12.648 27.856 13.392 ;
  LAYER M1 ;
        RECT 27.824 13.488 27.856 13.728 ;
  LAYER M1 ;
        RECT 27.824 13.824 27.856 14.568 ;
  LAYER M1 ;
        RECT 27.824 14.664 27.856 14.904 ;
  LAYER M1 ;
        RECT 27.824 15 27.856 15.744 ;
  LAYER M1 ;
        RECT 27.824 15.84 27.856 16.08 ;
  LAYER M1 ;
        RECT 27.824 16.176 27.856 16.92 ;
  LAYER M1 ;
        RECT 27.824 17.016 27.856 17.256 ;
  LAYER M1 ;
        RECT 27.824 17.352 27.856 18.096 ;
  LAYER M1 ;
        RECT 27.824 18.192 27.856 18.432 ;
  LAYER M1 ;
        RECT 27.824 18.528 27.856 19.272 ;
  LAYER M1 ;
        RECT 27.824 19.368 27.856 19.608 ;
  LAYER M1 ;
        RECT 27.824 19.704 27.856 20.448 ;
  LAYER M1 ;
        RECT 27.824 20.544 27.856 20.784 ;
  LAYER M1 ;
        RECT 27.824 20.88 27.856 21.624 ;
  LAYER M1 ;
        RECT 27.824 21.72 27.856 21.96 ;
  LAYER M1 ;
        RECT 27.824 22.056 27.856 22.8 ;
  LAYER M1 ;
        RECT 27.824 22.896 27.856 23.136 ;
  LAYER M1 ;
        RECT 27.824 23.232 27.856 23.976 ;
  LAYER M1 ;
        RECT 27.824 24.072 27.856 24.312 ;
  LAYER M1 ;
        RECT 27.824 24.576 27.856 24.816 ;
  LAYER M1 ;
        RECT 27.904 12.648 27.936 13.392 ;
  LAYER M1 ;
        RECT 27.904 13.824 27.936 14.568 ;
  LAYER M1 ;
        RECT 27.904 15 27.936 15.744 ;
  LAYER M1 ;
        RECT 27.904 16.176 27.936 16.92 ;
  LAYER M1 ;
        RECT 27.904 17.352 27.936 18.096 ;
  LAYER M1 ;
        RECT 27.904 18.528 27.936 19.272 ;
  LAYER M1 ;
        RECT 27.904 19.704 27.936 20.448 ;
  LAYER M1 ;
        RECT 27.904 20.88 27.936 21.624 ;
  LAYER M1 ;
        RECT 27.904 22.056 27.936 22.8 ;
  LAYER M1 ;
        RECT 27.904 23.232 27.936 23.976 ;
  LAYER M1 ;
        RECT 27.984 12.648 28.016 13.392 ;
  LAYER M1 ;
        RECT 27.984 13.488 28.016 13.728 ;
  LAYER M1 ;
        RECT 27.984 13.824 28.016 14.568 ;
  LAYER M1 ;
        RECT 27.984 14.664 28.016 14.904 ;
  LAYER M1 ;
        RECT 27.984 15 28.016 15.744 ;
  LAYER M1 ;
        RECT 27.984 15.84 28.016 16.08 ;
  LAYER M1 ;
        RECT 27.984 16.176 28.016 16.92 ;
  LAYER M1 ;
        RECT 27.984 17.016 28.016 17.256 ;
  LAYER M1 ;
        RECT 27.984 17.352 28.016 18.096 ;
  LAYER M1 ;
        RECT 27.984 18.192 28.016 18.432 ;
  LAYER M1 ;
        RECT 27.984 18.528 28.016 19.272 ;
  LAYER M1 ;
        RECT 27.984 19.368 28.016 19.608 ;
  LAYER M1 ;
        RECT 27.984 19.704 28.016 20.448 ;
  LAYER M1 ;
        RECT 27.984 20.544 28.016 20.784 ;
  LAYER M1 ;
        RECT 27.984 20.88 28.016 21.624 ;
  LAYER M1 ;
        RECT 27.984 21.72 28.016 21.96 ;
  LAYER M1 ;
        RECT 27.984 22.056 28.016 22.8 ;
  LAYER M1 ;
        RECT 27.984 22.896 28.016 23.136 ;
  LAYER M1 ;
        RECT 27.984 23.232 28.016 23.976 ;
  LAYER M1 ;
        RECT 27.984 24.072 28.016 24.312 ;
  LAYER M1 ;
        RECT 27.984 24.576 28.016 24.816 ;
  LAYER M1 ;
        RECT 28.064 12.648 28.096 13.392 ;
  LAYER M1 ;
        RECT 28.064 13.824 28.096 14.568 ;
  LAYER M1 ;
        RECT 28.064 15 28.096 15.744 ;
  LAYER M1 ;
        RECT 28.064 16.176 28.096 16.92 ;
  LAYER M1 ;
        RECT 28.064 17.352 28.096 18.096 ;
  LAYER M1 ;
        RECT 28.064 18.528 28.096 19.272 ;
  LAYER M1 ;
        RECT 28.064 19.704 28.096 20.448 ;
  LAYER M1 ;
        RECT 28.064 20.88 28.096 21.624 ;
  LAYER M1 ;
        RECT 28.064 22.056 28.096 22.8 ;
  LAYER M1 ;
        RECT 28.064 23.232 28.096 23.976 ;
  LAYER M1 ;
        RECT 28.144 12.648 28.176 13.392 ;
  LAYER M1 ;
        RECT 28.144 13.488 28.176 13.728 ;
  LAYER M1 ;
        RECT 28.144 13.824 28.176 14.568 ;
  LAYER M1 ;
        RECT 28.144 14.664 28.176 14.904 ;
  LAYER M1 ;
        RECT 28.144 15 28.176 15.744 ;
  LAYER M1 ;
        RECT 28.144 15.84 28.176 16.08 ;
  LAYER M1 ;
        RECT 28.144 16.176 28.176 16.92 ;
  LAYER M1 ;
        RECT 28.144 17.016 28.176 17.256 ;
  LAYER M1 ;
        RECT 28.144 17.352 28.176 18.096 ;
  LAYER M1 ;
        RECT 28.144 18.192 28.176 18.432 ;
  LAYER M1 ;
        RECT 28.144 18.528 28.176 19.272 ;
  LAYER M1 ;
        RECT 28.144 19.368 28.176 19.608 ;
  LAYER M1 ;
        RECT 28.144 19.704 28.176 20.448 ;
  LAYER M1 ;
        RECT 28.144 20.544 28.176 20.784 ;
  LAYER M1 ;
        RECT 28.144 20.88 28.176 21.624 ;
  LAYER M1 ;
        RECT 28.144 21.72 28.176 21.96 ;
  LAYER M1 ;
        RECT 28.144 22.056 28.176 22.8 ;
  LAYER M1 ;
        RECT 28.144 22.896 28.176 23.136 ;
  LAYER M1 ;
        RECT 28.144 23.232 28.176 23.976 ;
  LAYER M1 ;
        RECT 28.144 24.072 28.176 24.312 ;
  LAYER M1 ;
        RECT 28.144 24.576 28.176 24.816 ;
  LAYER M1 ;
        RECT 28.224 12.648 28.256 13.392 ;
  LAYER M1 ;
        RECT 28.224 13.824 28.256 14.568 ;
  LAYER M1 ;
        RECT 28.224 15 28.256 15.744 ;
  LAYER M1 ;
        RECT 28.224 16.176 28.256 16.92 ;
  LAYER M1 ;
        RECT 28.224 17.352 28.256 18.096 ;
  LAYER M1 ;
        RECT 28.224 18.528 28.256 19.272 ;
  LAYER M1 ;
        RECT 28.224 19.704 28.256 20.448 ;
  LAYER M1 ;
        RECT 28.224 20.88 28.256 21.624 ;
  LAYER M1 ;
        RECT 28.224 22.056 28.256 22.8 ;
  LAYER M1 ;
        RECT 28.224 23.232 28.256 23.976 ;
  LAYER M1 ;
        RECT 28.304 12.648 28.336 13.392 ;
  LAYER M1 ;
        RECT 28.304 13.488 28.336 13.728 ;
  LAYER M1 ;
        RECT 28.304 13.824 28.336 14.568 ;
  LAYER M1 ;
        RECT 28.304 14.664 28.336 14.904 ;
  LAYER M1 ;
        RECT 28.304 15 28.336 15.744 ;
  LAYER M1 ;
        RECT 28.304 15.84 28.336 16.08 ;
  LAYER M1 ;
        RECT 28.304 16.176 28.336 16.92 ;
  LAYER M1 ;
        RECT 28.304 17.016 28.336 17.256 ;
  LAYER M1 ;
        RECT 28.304 17.352 28.336 18.096 ;
  LAYER M1 ;
        RECT 28.304 18.192 28.336 18.432 ;
  LAYER M1 ;
        RECT 28.304 18.528 28.336 19.272 ;
  LAYER M1 ;
        RECT 28.304 19.368 28.336 19.608 ;
  LAYER M1 ;
        RECT 28.304 19.704 28.336 20.448 ;
  LAYER M1 ;
        RECT 28.304 20.544 28.336 20.784 ;
  LAYER M1 ;
        RECT 28.304 20.88 28.336 21.624 ;
  LAYER M1 ;
        RECT 28.304 21.72 28.336 21.96 ;
  LAYER M1 ;
        RECT 28.304 22.056 28.336 22.8 ;
  LAYER M1 ;
        RECT 28.304 22.896 28.336 23.136 ;
  LAYER M1 ;
        RECT 28.304 23.232 28.336 23.976 ;
  LAYER M1 ;
        RECT 28.304 24.072 28.336 24.312 ;
  LAYER M1 ;
        RECT 28.304 24.576 28.336 24.816 ;
  LAYER M1 ;
        RECT 28.384 12.648 28.416 13.392 ;
  LAYER M1 ;
        RECT 28.384 13.824 28.416 14.568 ;
  LAYER M1 ;
        RECT 28.384 15 28.416 15.744 ;
  LAYER M1 ;
        RECT 28.384 16.176 28.416 16.92 ;
  LAYER M1 ;
        RECT 28.384 17.352 28.416 18.096 ;
  LAYER M1 ;
        RECT 28.384 18.528 28.416 19.272 ;
  LAYER M1 ;
        RECT 28.384 19.704 28.416 20.448 ;
  LAYER M1 ;
        RECT 28.384 20.88 28.416 21.624 ;
  LAYER M1 ;
        RECT 28.384 22.056 28.416 22.8 ;
  LAYER M1 ;
        RECT 28.384 23.232 28.416 23.976 ;
  LAYER M1 ;
        RECT 28.464 12.648 28.496 13.392 ;
  LAYER M1 ;
        RECT 28.464 13.488 28.496 13.728 ;
  LAYER M1 ;
        RECT 28.464 13.824 28.496 14.568 ;
  LAYER M1 ;
        RECT 28.464 14.664 28.496 14.904 ;
  LAYER M1 ;
        RECT 28.464 15 28.496 15.744 ;
  LAYER M1 ;
        RECT 28.464 15.84 28.496 16.08 ;
  LAYER M1 ;
        RECT 28.464 16.176 28.496 16.92 ;
  LAYER M1 ;
        RECT 28.464 17.016 28.496 17.256 ;
  LAYER M1 ;
        RECT 28.464 17.352 28.496 18.096 ;
  LAYER M1 ;
        RECT 28.464 18.192 28.496 18.432 ;
  LAYER M1 ;
        RECT 28.464 18.528 28.496 19.272 ;
  LAYER M1 ;
        RECT 28.464 19.368 28.496 19.608 ;
  LAYER M1 ;
        RECT 28.464 19.704 28.496 20.448 ;
  LAYER M1 ;
        RECT 28.464 20.544 28.496 20.784 ;
  LAYER M1 ;
        RECT 28.464 20.88 28.496 21.624 ;
  LAYER M1 ;
        RECT 28.464 21.72 28.496 21.96 ;
  LAYER M1 ;
        RECT 28.464 22.056 28.496 22.8 ;
  LAYER M1 ;
        RECT 28.464 22.896 28.496 23.136 ;
  LAYER M1 ;
        RECT 28.464 23.232 28.496 23.976 ;
  LAYER M1 ;
        RECT 28.464 24.072 28.496 24.312 ;
  LAYER M1 ;
        RECT 28.464 24.576 28.496 24.816 ;
  LAYER M1 ;
        RECT 28.544 12.648 28.576 13.392 ;
  LAYER M1 ;
        RECT 28.544 13.824 28.576 14.568 ;
  LAYER M1 ;
        RECT 28.544 15 28.576 15.744 ;
  LAYER M1 ;
        RECT 28.544 16.176 28.576 16.92 ;
  LAYER M1 ;
        RECT 28.544 17.352 28.576 18.096 ;
  LAYER M1 ;
        RECT 28.544 18.528 28.576 19.272 ;
  LAYER M1 ;
        RECT 28.544 19.704 28.576 20.448 ;
  LAYER M1 ;
        RECT 28.544 20.88 28.576 21.624 ;
  LAYER M1 ;
        RECT 28.544 22.056 28.576 22.8 ;
  LAYER M1 ;
        RECT 28.544 23.232 28.576 23.976 ;
  LAYER M1 ;
        RECT 28.624 12.648 28.656 13.392 ;
  LAYER M1 ;
        RECT 28.624 13.488 28.656 13.728 ;
  LAYER M1 ;
        RECT 28.624 13.824 28.656 14.568 ;
  LAYER M1 ;
        RECT 28.624 14.664 28.656 14.904 ;
  LAYER M1 ;
        RECT 28.624 15 28.656 15.744 ;
  LAYER M1 ;
        RECT 28.624 15.84 28.656 16.08 ;
  LAYER M1 ;
        RECT 28.624 16.176 28.656 16.92 ;
  LAYER M1 ;
        RECT 28.624 17.016 28.656 17.256 ;
  LAYER M1 ;
        RECT 28.624 17.352 28.656 18.096 ;
  LAYER M1 ;
        RECT 28.624 18.192 28.656 18.432 ;
  LAYER M1 ;
        RECT 28.624 18.528 28.656 19.272 ;
  LAYER M1 ;
        RECT 28.624 19.368 28.656 19.608 ;
  LAYER M1 ;
        RECT 28.624 19.704 28.656 20.448 ;
  LAYER M1 ;
        RECT 28.624 20.544 28.656 20.784 ;
  LAYER M1 ;
        RECT 28.624 20.88 28.656 21.624 ;
  LAYER M1 ;
        RECT 28.624 21.72 28.656 21.96 ;
  LAYER M1 ;
        RECT 28.624 22.056 28.656 22.8 ;
  LAYER M1 ;
        RECT 28.624 22.896 28.656 23.136 ;
  LAYER M1 ;
        RECT 28.624 23.232 28.656 23.976 ;
  LAYER M1 ;
        RECT 28.624 24.072 28.656 24.312 ;
  LAYER M1 ;
        RECT 28.624 24.576 28.656 24.816 ;
  LAYER M1 ;
        RECT 28.704 12.648 28.736 13.392 ;
  LAYER M1 ;
        RECT 28.704 13.824 28.736 14.568 ;
  LAYER M1 ;
        RECT 28.704 15 28.736 15.744 ;
  LAYER M1 ;
        RECT 28.704 16.176 28.736 16.92 ;
  LAYER M1 ;
        RECT 28.704 17.352 28.736 18.096 ;
  LAYER M1 ;
        RECT 28.704 18.528 28.736 19.272 ;
  LAYER M1 ;
        RECT 28.704 19.704 28.736 20.448 ;
  LAYER M1 ;
        RECT 28.704 20.88 28.736 21.624 ;
  LAYER M1 ;
        RECT 28.704 22.056 28.736 22.8 ;
  LAYER M1 ;
        RECT 28.704 23.232 28.736 23.976 ;
  LAYER M1 ;
        RECT 28.784 12.648 28.816 13.392 ;
  LAYER M1 ;
        RECT 28.784 13.488 28.816 13.728 ;
  LAYER M1 ;
        RECT 28.784 13.824 28.816 14.568 ;
  LAYER M1 ;
        RECT 28.784 14.664 28.816 14.904 ;
  LAYER M1 ;
        RECT 28.784 15 28.816 15.744 ;
  LAYER M1 ;
        RECT 28.784 15.84 28.816 16.08 ;
  LAYER M1 ;
        RECT 28.784 16.176 28.816 16.92 ;
  LAYER M1 ;
        RECT 28.784 17.016 28.816 17.256 ;
  LAYER M1 ;
        RECT 28.784 17.352 28.816 18.096 ;
  LAYER M1 ;
        RECT 28.784 18.192 28.816 18.432 ;
  LAYER M1 ;
        RECT 28.784 18.528 28.816 19.272 ;
  LAYER M1 ;
        RECT 28.784 19.368 28.816 19.608 ;
  LAYER M1 ;
        RECT 28.784 19.704 28.816 20.448 ;
  LAYER M1 ;
        RECT 28.784 20.544 28.816 20.784 ;
  LAYER M1 ;
        RECT 28.784 20.88 28.816 21.624 ;
  LAYER M1 ;
        RECT 28.784 21.72 28.816 21.96 ;
  LAYER M1 ;
        RECT 28.784 22.056 28.816 22.8 ;
  LAYER M1 ;
        RECT 28.784 22.896 28.816 23.136 ;
  LAYER M1 ;
        RECT 28.784 23.232 28.816 23.976 ;
  LAYER M1 ;
        RECT 28.784 24.072 28.816 24.312 ;
  LAYER M1 ;
        RECT 28.784 24.576 28.816 24.816 ;
  LAYER M1 ;
        RECT 28.864 12.648 28.896 13.392 ;
  LAYER M1 ;
        RECT 28.864 13.824 28.896 14.568 ;
  LAYER M1 ;
        RECT 28.864 15 28.896 15.744 ;
  LAYER M1 ;
        RECT 28.864 16.176 28.896 16.92 ;
  LAYER M1 ;
        RECT 28.864 17.352 28.896 18.096 ;
  LAYER M1 ;
        RECT 28.864 18.528 28.896 19.272 ;
  LAYER M1 ;
        RECT 28.864 19.704 28.896 20.448 ;
  LAYER M1 ;
        RECT 28.864 20.88 28.896 21.624 ;
  LAYER M1 ;
        RECT 28.864 22.056 28.896 22.8 ;
  LAYER M1 ;
        RECT 28.864 23.232 28.896 23.976 ;
  LAYER M1 ;
        RECT 28.944 12.648 28.976 13.392 ;
  LAYER M1 ;
        RECT 28.944 13.488 28.976 13.728 ;
  LAYER M1 ;
        RECT 28.944 13.824 28.976 14.568 ;
  LAYER M1 ;
        RECT 28.944 14.664 28.976 14.904 ;
  LAYER M1 ;
        RECT 28.944 15 28.976 15.744 ;
  LAYER M1 ;
        RECT 28.944 15.84 28.976 16.08 ;
  LAYER M1 ;
        RECT 28.944 16.176 28.976 16.92 ;
  LAYER M1 ;
        RECT 28.944 17.016 28.976 17.256 ;
  LAYER M1 ;
        RECT 28.944 17.352 28.976 18.096 ;
  LAYER M1 ;
        RECT 28.944 18.192 28.976 18.432 ;
  LAYER M1 ;
        RECT 28.944 18.528 28.976 19.272 ;
  LAYER M1 ;
        RECT 28.944 19.368 28.976 19.608 ;
  LAYER M1 ;
        RECT 28.944 19.704 28.976 20.448 ;
  LAYER M1 ;
        RECT 28.944 20.544 28.976 20.784 ;
  LAYER M1 ;
        RECT 28.944 20.88 28.976 21.624 ;
  LAYER M1 ;
        RECT 28.944 21.72 28.976 21.96 ;
  LAYER M1 ;
        RECT 28.944 22.056 28.976 22.8 ;
  LAYER M1 ;
        RECT 28.944 22.896 28.976 23.136 ;
  LAYER M1 ;
        RECT 28.944 23.232 28.976 23.976 ;
  LAYER M1 ;
        RECT 28.944 24.072 28.976 24.312 ;
  LAYER M1 ;
        RECT 28.944 24.576 28.976 24.816 ;
  LAYER M1 ;
        RECT 29.024 12.648 29.056 13.392 ;
  LAYER M1 ;
        RECT 29.024 13.824 29.056 14.568 ;
  LAYER M1 ;
        RECT 29.024 15 29.056 15.744 ;
  LAYER M1 ;
        RECT 29.024 16.176 29.056 16.92 ;
  LAYER M1 ;
        RECT 29.024 17.352 29.056 18.096 ;
  LAYER M1 ;
        RECT 29.024 18.528 29.056 19.272 ;
  LAYER M1 ;
        RECT 29.024 19.704 29.056 20.448 ;
  LAYER M1 ;
        RECT 29.024 20.88 29.056 21.624 ;
  LAYER M1 ;
        RECT 29.024 22.056 29.056 22.8 ;
  LAYER M1 ;
        RECT 29.024 23.232 29.056 23.976 ;
  LAYER M1 ;
        RECT 29.104 12.648 29.136 13.392 ;
  LAYER M1 ;
        RECT 29.104 13.488 29.136 13.728 ;
  LAYER M1 ;
        RECT 29.104 13.824 29.136 14.568 ;
  LAYER M1 ;
        RECT 29.104 14.664 29.136 14.904 ;
  LAYER M1 ;
        RECT 29.104 15 29.136 15.744 ;
  LAYER M1 ;
        RECT 29.104 15.84 29.136 16.08 ;
  LAYER M1 ;
        RECT 29.104 16.176 29.136 16.92 ;
  LAYER M1 ;
        RECT 29.104 17.016 29.136 17.256 ;
  LAYER M1 ;
        RECT 29.104 17.352 29.136 18.096 ;
  LAYER M1 ;
        RECT 29.104 18.192 29.136 18.432 ;
  LAYER M1 ;
        RECT 29.104 18.528 29.136 19.272 ;
  LAYER M1 ;
        RECT 29.104 19.368 29.136 19.608 ;
  LAYER M1 ;
        RECT 29.104 19.704 29.136 20.448 ;
  LAYER M1 ;
        RECT 29.104 20.544 29.136 20.784 ;
  LAYER M1 ;
        RECT 29.104 20.88 29.136 21.624 ;
  LAYER M1 ;
        RECT 29.104 21.72 29.136 21.96 ;
  LAYER M1 ;
        RECT 29.104 22.056 29.136 22.8 ;
  LAYER M1 ;
        RECT 29.104 22.896 29.136 23.136 ;
  LAYER M1 ;
        RECT 29.104 23.232 29.136 23.976 ;
  LAYER M1 ;
        RECT 29.104 24.072 29.136 24.312 ;
  LAYER M1 ;
        RECT 29.104 24.576 29.136 24.816 ;
  LAYER M1 ;
        RECT 29.184 12.648 29.216 13.392 ;
  LAYER M1 ;
        RECT 29.184 13.824 29.216 14.568 ;
  LAYER M1 ;
        RECT 29.184 15 29.216 15.744 ;
  LAYER M1 ;
        RECT 29.184 16.176 29.216 16.92 ;
  LAYER M1 ;
        RECT 29.184 17.352 29.216 18.096 ;
  LAYER M1 ;
        RECT 29.184 18.528 29.216 19.272 ;
  LAYER M1 ;
        RECT 29.184 19.704 29.216 20.448 ;
  LAYER M1 ;
        RECT 29.184 20.88 29.216 21.624 ;
  LAYER M1 ;
        RECT 29.184 22.056 29.216 22.8 ;
  LAYER M1 ;
        RECT 29.184 23.232 29.216 23.976 ;
  LAYER M1 ;
        RECT 29.264 12.648 29.296 13.392 ;
  LAYER M1 ;
        RECT 29.264 13.488 29.296 13.728 ;
  LAYER M1 ;
        RECT 29.264 13.824 29.296 14.568 ;
  LAYER M1 ;
        RECT 29.264 14.664 29.296 14.904 ;
  LAYER M1 ;
        RECT 29.264 15 29.296 15.744 ;
  LAYER M1 ;
        RECT 29.264 15.84 29.296 16.08 ;
  LAYER M1 ;
        RECT 29.264 16.176 29.296 16.92 ;
  LAYER M1 ;
        RECT 29.264 17.016 29.296 17.256 ;
  LAYER M1 ;
        RECT 29.264 17.352 29.296 18.096 ;
  LAYER M1 ;
        RECT 29.264 18.192 29.296 18.432 ;
  LAYER M1 ;
        RECT 29.264 18.528 29.296 19.272 ;
  LAYER M1 ;
        RECT 29.264 19.368 29.296 19.608 ;
  LAYER M1 ;
        RECT 29.264 19.704 29.296 20.448 ;
  LAYER M1 ;
        RECT 29.264 20.544 29.296 20.784 ;
  LAYER M1 ;
        RECT 29.264 20.88 29.296 21.624 ;
  LAYER M1 ;
        RECT 29.264 21.72 29.296 21.96 ;
  LAYER M1 ;
        RECT 29.264 22.056 29.296 22.8 ;
  LAYER M1 ;
        RECT 29.264 22.896 29.296 23.136 ;
  LAYER M1 ;
        RECT 29.264 23.232 29.296 23.976 ;
  LAYER M1 ;
        RECT 29.264 24.072 29.296 24.312 ;
  LAYER M1 ;
        RECT 29.264 24.576 29.296 24.816 ;
  LAYER M1 ;
        RECT 29.344 12.648 29.376 13.392 ;
  LAYER M1 ;
        RECT 29.344 13.824 29.376 14.568 ;
  LAYER M1 ;
        RECT 29.344 15 29.376 15.744 ;
  LAYER M1 ;
        RECT 29.344 16.176 29.376 16.92 ;
  LAYER M1 ;
        RECT 29.344 17.352 29.376 18.096 ;
  LAYER M1 ;
        RECT 29.344 18.528 29.376 19.272 ;
  LAYER M1 ;
        RECT 29.344 19.704 29.376 20.448 ;
  LAYER M1 ;
        RECT 29.344 20.88 29.376 21.624 ;
  LAYER M1 ;
        RECT 29.344 22.056 29.376 22.8 ;
  LAYER M1 ;
        RECT 29.344 23.232 29.376 23.976 ;
  LAYER M1 ;
        RECT 29.424 12.648 29.456 13.392 ;
  LAYER M1 ;
        RECT 29.424 13.488 29.456 13.728 ;
  LAYER M1 ;
        RECT 29.424 13.824 29.456 14.568 ;
  LAYER M1 ;
        RECT 29.424 14.664 29.456 14.904 ;
  LAYER M1 ;
        RECT 29.424 15 29.456 15.744 ;
  LAYER M1 ;
        RECT 29.424 15.84 29.456 16.08 ;
  LAYER M1 ;
        RECT 29.424 16.176 29.456 16.92 ;
  LAYER M1 ;
        RECT 29.424 17.016 29.456 17.256 ;
  LAYER M1 ;
        RECT 29.424 17.352 29.456 18.096 ;
  LAYER M1 ;
        RECT 29.424 18.192 29.456 18.432 ;
  LAYER M1 ;
        RECT 29.424 18.528 29.456 19.272 ;
  LAYER M1 ;
        RECT 29.424 19.368 29.456 19.608 ;
  LAYER M1 ;
        RECT 29.424 19.704 29.456 20.448 ;
  LAYER M1 ;
        RECT 29.424 20.544 29.456 20.784 ;
  LAYER M1 ;
        RECT 29.424 20.88 29.456 21.624 ;
  LAYER M1 ;
        RECT 29.424 21.72 29.456 21.96 ;
  LAYER M1 ;
        RECT 29.424 22.056 29.456 22.8 ;
  LAYER M1 ;
        RECT 29.424 22.896 29.456 23.136 ;
  LAYER M1 ;
        RECT 29.424 23.232 29.456 23.976 ;
  LAYER M1 ;
        RECT 29.424 24.072 29.456 24.312 ;
  LAYER M1 ;
        RECT 29.424 24.576 29.456 24.816 ;
  LAYER M1 ;
        RECT 29.504 12.648 29.536 13.392 ;
  LAYER M1 ;
        RECT 29.504 13.824 29.536 14.568 ;
  LAYER M1 ;
        RECT 29.504 15 29.536 15.744 ;
  LAYER M1 ;
        RECT 29.504 16.176 29.536 16.92 ;
  LAYER M1 ;
        RECT 29.504 17.352 29.536 18.096 ;
  LAYER M1 ;
        RECT 29.504 18.528 29.536 19.272 ;
  LAYER M1 ;
        RECT 29.504 19.704 29.536 20.448 ;
  LAYER M1 ;
        RECT 29.504 20.88 29.536 21.624 ;
  LAYER M1 ;
        RECT 29.504 22.056 29.536 22.8 ;
  LAYER M1 ;
        RECT 29.504 23.232 29.536 23.976 ;
  LAYER M1 ;
        RECT 29.584 12.648 29.616 13.392 ;
  LAYER M1 ;
        RECT 29.584 13.488 29.616 13.728 ;
  LAYER M1 ;
        RECT 29.584 13.824 29.616 14.568 ;
  LAYER M1 ;
        RECT 29.584 14.664 29.616 14.904 ;
  LAYER M1 ;
        RECT 29.584 15 29.616 15.744 ;
  LAYER M1 ;
        RECT 29.584 15.84 29.616 16.08 ;
  LAYER M1 ;
        RECT 29.584 16.176 29.616 16.92 ;
  LAYER M1 ;
        RECT 29.584 17.016 29.616 17.256 ;
  LAYER M1 ;
        RECT 29.584 17.352 29.616 18.096 ;
  LAYER M1 ;
        RECT 29.584 18.192 29.616 18.432 ;
  LAYER M1 ;
        RECT 29.584 18.528 29.616 19.272 ;
  LAYER M1 ;
        RECT 29.584 19.368 29.616 19.608 ;
  LAYER M1 ;
        RECT 29.584 19.704 29.616 20.448 ;
  LAYER M1 ;
        RECT 29.584 20.544 29.616 20.784 ;
  LAYER M1 ;
        RECT 29.584 20.88 29.616 21.624 ;
  LAYER M1 ;
        RECT 29.584 21.72 29.616 21.96 ;
  LAYER M1 ;
        RECT 29.584 22.056 29.616 22.8 ;
  LAYER M1 ;
        RECT 29.584 22.896 29.616 23.136 ;
  LAYER M1 ;
        RECT 29.584 23.232 29.616 23.976 ;
  LAYER M1 ;
        RECT 29.584 24.072 29.616 24.312 ;
  LAYER M1 ;
        RECT 29.584 24.576 29.616 24.816 ;
  LAYER M1 ;
        RECT 29.664 12.648 29.696 13.392 ;
  LAYER M1 ;
        RECT 29.664 13.824 29.696 14.568 ;
  LAYER M1 ;
        RECT 29.664 15 29.696 15.744 ;
  LAYER M1 ;
        RECT 29.664 16.176 29.696 16.92 ;
  LAYER M1 ;
        RECT 29.664 17.352 29.696 18.096 ;
  LAYER M1 ;
        RECT 29.664 18.528 29.696 19.272 ;
  LAYER M1 ;
        RECT 29.664 19.704 29.696 20.448 ;
  LAYER M1 ;
        RECT 29.664 20.88 29.696 21.624 ;
  LAYER M1 ;
        RECT 29.664 22.056 29.696 22.8 ;
  LAYER M1 ;
        RECT 29.664 23.232 29.696 23.976 ;
  LAYER M1 ;
        RECT 29.744 12.648 29.776 13.392 ;
  LAYER M1 ;
        RECT 29.744 13.488 29.776 13.728 ;
  LAYER M1 ;
        RECT 29.744 13.824 29.776 14.568 ;
  LAYER M1 ;
        RECT 29.744 14.664 29.776 14.904 ;
  LAYER M1 ;
        RECT 29.744 15 29.776 15.744 ;
  LAYER M1 ;
        RECT 29.744 15.84 29.776 16.08 ;
  LAYER M1 ;
        RECT 29.744 16.176 29.776 16.92 ;
  LAYER M1 ;
        RECT 29.744 17.016 29.776 17.256 ;
  LAYER M1 ;
        RECT 29.744 17.352 29.776 18.096 ;
  LAYER M1 ;
        RECT 29.744 18.192 29.776 18.432 ;
  LAYER M1 ;
        RECT 29.744 18.528 29.776 19.272 ;
  LAYER M1 ;
        RECT 29.744 19.368 29.776 19.608 ;
  LAYER M1 ;
        RECT 29.744 19.704 29.776 20.448 ;
  LAYER M1 ;
        RECT 29.744 20.544 29.776 20.784 ;
  LAYER M1 ;
        RECT 29.744 20.88 29.776 21.624 ;
  LAYER M1 ;
        RECT 29.744 21.72 29.776 21.96 ;
  LAYER M1 ;
        RECT 29.744 22.056 29.776 22.8 ;
  LAYER M1 ;
        RECT 29.744 22.896 29.776 23.136 ;
  LAYER M1 ;
        RECT 29.744 23.232 29.776 23.976 ;
  LAYER M1 ;
        RECT 29.744 24.072 29.776 24.312 ;
  LAYER M1 ;
        RECT 29.744 24.576 29.776 24.816 ;
  LAYER M1 ;
        RECT 29.824 12.648 29.856 13.392 ;
  LAYER M1 ;
        RECT 29.824 13.824 29.856 14.568 ;
  LAYER M1 ;
        RECT 29.824 15 29.856 15.744 ;
  LAYER M1 ;
        RECT 29.824 16.176 29.856 16.92 ;
  LAYER M1 ;
        RECT 29.824 17.352 29.856 18.096 ;
  LAYER M1 ;
        RECT 29.824 18.528 29.856 19.272 ;
  LAYER M1 ;
        RECT 29.824 19.704 29.856 20.448 ;
  LAYER M1 ;
        RECT 29.824 20.88 29.856 21.624 ;
  LAYER M1 ;
        RECT 29.824 22.056 29.856 22.8 ;
  LAYER M1 ;
        RECT 29.824 23.232 29.856 23.976 ;
  LAYER M1 ;
        RECT 29.904 12.648 29.936 13.392 ;
  LAYER M1 ;
        RECT 29.904 13.488 29.936 13.728 ;
  LAYER M1 ;
        RECT 29.904 13.824 29.936 14.568 ;
  LAYER M1 ;
        RECT 29.904 14.664 29.936 14.904 ;
  LAYER M1 ;
        RECT 29.904 15 29.936 15.744 ;
  LAYER M1 ;
        RECT 29.904 15.84 29.936 16.08 ;
  LAYER M1 ;
        RECT 29.904 16.176 29.936 16.92 ;
  LAYER M1 ;
        RECT 29.904 17.016 29.936 17.256 ;
  LAYER M1 ;
        RECT 29.904 17.352 29.936 18.096 ;
  LAYER M1 ;
        RECT 29.904 18.192 29.936 18.432 ;
  LAYER M1 ;
        RECT 29.904 18.528 29.936 19.272 ;
  LAYER M1 ;
        RECT 29.904 19.368 29.936 19.608 ;
  LAYER M1 ;
        RECT 29.904 19.704 29.936 20.448 ;
  LAYER M1 ;
        RECT 29.904 20.544 29.936 20.784 ;
  LAYER M1 ;
        RECT 29.904 20.88 29.936 21.624 ;
  LAYER M1 ;
        RECT 29.904 21.72 29.936 21.96 ;
  LAYER M1 ;
        RECT 29.904 22.056 29.936 22.8 ;
  LAYER M1 ;
        RECT 29.904 22.896 29.936 23.136 ;
  LAYER M1 ;
        RECT 29.904 23.232 29.936 23.976 ;
  LAYER M1 ;
        RECT 29.904 24.072 29.936 24.312 ;
  LAYER M1 ;
        RECT 29.904 24.576 29.936 24.816 ;
  LAYER M1 ;
        RECT 29.984 12.648 30.016 13.392 ;
  LAYER M1 ;
        RECT 29.984 13.824 30.016 14.568 ;
  LAYER M1 ;
        RECT 29.984 15 30.016 15.744 ;
  LAYER M1 ;
        RECT 29.984 16.176 30.016 16.92 ;
  LAYER M1 ;
        RECT 29.984 17.352 30.016 18.096 ;
  LAYER M1 ;
        RECT 29.984 18.528 30.016 19.272 ;
  LAYER M1 ;
        RECT 29.984 19.704 30.016 20.448 ;
  LAYER M1 ;
        RECT 29.984 20.88 30.016 21.624 ;
  LAYER M1 ;
        RECT 29.984 22.056 30.016 22.8 ;
  LAYER M1 ;
        RECT 29.984 23.232 30.016 23.976 ;
  LAYER M1 ;
        RECT 30.064 12.648 30.096 13.392 ;
  LAYER M1 ;
        RECT 30.064 13.488 30.096 13.728 ;
  LAYER M1 ;
        RECT 30.064 13.824 30.096 14.568 ;
  LAYER M1 ;
        RECT 30.064 14.664 30.096 14.904 ;
  LAYER M1 ;
        RECT 30.064 15 30.096 15.744 ;
  LAYER M1 ;
        RECT 30.064 15.84 30.096 16.08 ;
  LAYER M1 ;
        RECT 30.064 16.176 30.096 16.92 ;
  LAYER M1 ;
        RECT 30.064 17.016 30.096 17.256 ;
  LAYER M1 ;
        RECT 30.064 17.352 30.096 18.096 ;
  LAYER M1 ;
        RECT 30.064 18.192 30.096 18.432 ;
  LAYER M1 ;
        RECT 30.064 18.528 30.096 19.272 ;
  LAYER M1 ;
        RECT 30.064 19.368 30.096 19.608 ;
  LAYER M1 ;
        RECT 30.064 19.704 30.096 20.448 ;
  LAYER M1 ;
        RECT 30.064 20.544 30.096 20.784 ;
  LAYER M1 ;
        RECT 30.064 20.88 30.096 21.624 ;
  LAYER M1 ;
        RECT 30.064 21.72 30.096 21.96 ;
  LAYER M1 ;
        RECT 30.064 22.056 30.096 22.8 ;
  LAYER M1 ;
        RECT 30.064 22.896 30.096 23.136 ;
  LAYER M1 ;
        RECT 30.064 23.232 30.096 23.976 ;
  LAYER M1 ;
        RECT 30.064 24.072 30.096 24.312 ;
  LAYER M1 ;
        RECT 30.064 24.576 30.096 24.816 ;
  LAYER M1 ;
        RECT 30.144 12.648 30.176 13.392 ;
  LAYER M1 ;
        RECT 30.144 13.824 30.176 14.568 ;
  LAYER M1 ;
        RECT 30.144 15 30.176 15.744 ;
  LAYER M1 ;
        RECT 30.144 16.176 30.176 16.92 ;
  LAYER M1 ;
        RECT 30.144 17.352 30.176 18.096 ;
  LAYER M1 ;
        RECT 30.144 18.528 30.176 19.272 ;
  LAYER M1 ;
        RECT 30.144 19.704 30.176 20.448 ;
  LAYER M1 ;
        RECT 30.144 20.88 30.176 21.624 ;
  LAYER M1 ;
        RECT 30.144 22.056 30.176 22.8 ;
  LAYER M1 ;
        RECT 30.144 23.232 30.176 23.976 ;
  LAYER M1 ;
        RECT 30.224 12.648 30.256 13.392 ;
  LAYER M1 ;
        RECT 30.224 13.488 30.256 13.728 ;
  LAYER M1 ;
        RECT 30.224 13.824 30.256 14.568 ;
  LAYER M1 ;
        RECT 30.224 14.664 30.256 14.904 ;
  LAYER M1 ;
        RECT 30.224 15 30.256 15.744 ;
  LAYER M1 ;
        RECT 30.224 15.84 30.256 16.08 ;
  LAYER M1 ;
        RECT 30.224 16.176 30.256 16.92 ;
  LAYER M1 ;
        RECT 30.224 17.016 30.256 17.256 ;
  LAYER M1 ;
        RECT 30.224 17.352 30.256 18.096 ;
  LAYER M1 ;
        RECT 30.224 18.192 30.256 18.432 ;
  LAYER M1 ;
        RECT 30.224 18.528 30.256 19.272 ;
  LAYER M1 ;
        RECT 30.224 19.368 30.256 19.608 ;
  LAYER M1 ;
        RECT 30.224 19.704 30.256 20.448 ;
  LAYER M1 ;
        RECT 30.224 20.544 30.256 20.784 ;
  LAYER M1 ;
        RECT 30.224 20.88 30.256 21.624 ;
  LAYER M1 ;
        RECT 30.224 21.72 30.256 21.96 ;
  LAYER M1 ;
        RECT 30.224 22.056 30.256 22.8 ;
  LAYER M1 ;
        RECT 30.224 22.896 30.256 23.136 ;
  LAYER M1 ;
        RECT 30.224 23.232 30.256 23.976 ;
  LAYER M1 ;
        RECT 30.224 24.072 30.256 24.312 ;
  LAYER M1 ;
        RECT 30.224 24.576 30.256 24.816 ;
  LAYER M1 ;
        RECT 30.304 12.648 30.336 13.392 ;
  LAYER M1 ;
        RECT 30.304 13.824 30.336 14.568 ;
  LAYER M1 ;
        RECT 30.304 15 30.336 15.744 ;
  LAYER M1 ;
        RECT 30.304 16.176 30.336 16.92 ;
  LAYER M1 ;
        RECT 30.304 17.352 30.336 18.096 ;
  LAYER M1 ;
        RECT 30.304 18.528 30.336 19.272 ;
  LAYER M1 ;
        RECT 30.304 19.704 30.336 20.448 ;
  LAYER M1 ;
        RECT 30.304 20.88 30.336 21.624 ;
  LAYER M1 ;
        RECT 30.304 22.056 30.336 22.8 ;
  LAYER M1 ;
        RECT 30.304 23.232 30.336 23.976 ;
  LAYER M1 ;
        RECT 30.384 12.648 30.416 13.392 ;
  LAYER M1 ;
        RECT 30.384 13.488 30.416 13.728 ;
  LAYER M1 ;
        RECT 30.384 13.824 30.416 14.568 ;
  LAYER M1 ;
        RECT 30.384 14.664 30.416 14.904 ;
  LAYER M1 ;
        RECT 30.384 15 30.416 15.744 ;
  LAYER M1 ;
        RECT 30.384 15.84 30.416 16.08 ;
  LAYER M1 ;
        RECT 30.384 16.176 30.416 16.92 ;
  LAYER M1 ;
        RECT 30.384 17.016 30.416 17.256 ;
  LAYER M1 ;
        RECT 30.384 17.352 30.416 18.096 ;
  LAYER M1 ;
        RECT 30.384 18.192 30.416 18.432 ;
  LAYER M1 ;
        RECT 30.384 18.528 30.416 19.272 ;
  LAYER M1 ;
        RECT 30.384 19.368 30.416 19.608 ;
  LAYER M1 ;
        RECT 30.384 19.704 30.416 20.448 ;
  LAYER M1 ;
        RECT 30.384 20.544 30.416 20.784 ;
  LAYER M1 ;
        RECT 30.384 20.88 30.416 21.624 ;
  LAYER M1 ;
        RECT 30.384 21.72 30.416 21.96 ;
  LAYER M1 ;
        RECT 30.384 22.056 30.416 22.8 ;
  LAYER M1 ;
        RECT 30.384 22.896 30.416 23.136 ;
  LAYER M1 ;
        RECT 30.384 23.232 30.416 23.976 ;
  LAYER M1 ;
        RECT 30.384 24.072 30.416 24.312 ;
  LAYER M1 ;
        RECT 30.384 24.576 30.416 24.816 ;
  LAYER M1 ;
        RECT 30.464 12.648 30.496 13.392 ;
  LAYER M1 ;
        RECT 30.464 13.824 30.496 14.568 ;
  LAYER M1 ;
        RECT 30.464 15 30.496 15.744 ;
  LAYER M1 ;
        RECT 30.464 16.176 30.496 16.92 ;
  LAYER M1 ;
        RECT 30.464 17.352 30.496 18.096 ;
  LAYER M1 ;
        RECT 30.464 18.528 30.496 19.272 ;
  LAYER M1 ;
        RECT 30.464 19.704 30.496 20.448 ;
  LAYER M1 ;
        RECT 30.464 20.88 30.496 21.624 ;
  LAYER M1 ;
        RECT 30.464 22.056 30.496 22.8 ;
  LAYER M1 ;
        RECT 30.464 23.232 30.496 23.976 ;
  LAYER M1 ;
        RECT 30.544 12.648 30.576 13.392 ;
  LAYER M1 ;
        RECT 30.544 13.488 30.576 13.728 ;
  LAYER M1 ;
        RECT 30.544 13.824 30.576 14.568 ;
  LAYER M1 ;
        RECT 30.544 14.664 30.576 14.904 ;
  LAYER M1 ;
        RECT 30.544 15 30.576 15.744 ;
  LAYER M1 ;
        RECT 30.544 15.84 30.576 16.08 ;
  LAYER M1 ;
        RECT 30.544 16.176 30.576 16.92 ;
  LAYER M1 ;
        RECT 30.544 17.016 30.576 17.256 ;
  LAYER M1 ;
        RECT 30.544 17.352 30.576 18.096 ;
  LAYER M1 ;
        RECT 30.544 18.192 30.576 18.432 ;
  LAYER M1 ;
        RECT 30.544 18.528 30.576 19.272 ;
  LAYER M1 ;
        RECT 30.544 19.368 30.576 19.608 ;
  LAYER M1 ;
        RECT 30.544 19.704 30.576 20.448 ;
  LAYER M1 ;
        RECT 30.544 20.544 30.576 20.784 ;
  LAYER M1 ;
        RECT 30.544 20.88 30.576 21.624 ;
  LAYER M1 ;
        RECT 30.544 21.72 30.576 21.96 ;
  LAYER M1 ;
        RECT 30.544 22.056 30.576 22.8 ;
  LAYER M1 ;
        RECT 30.544 22.896 30.576 23.136 ;
  LAYER M1 ;
        RECT 30.544 23.232 30.576 23.976 ;
  LAYER M1 ;
        RECT 30.544 24.072 30.576 24.312 ;
  LAYER M1 ;
        RECT 30.544 24.576 30.576 24.816 ;
  LAYER M1 ;
        RECT 30.624 12.648 30.656 13.392 ;
  LAYER M1 ;
        RECT 30.624 13.824 30.656 14.568 ;
  LAYER M1 ;
        RECT 30.624 15 30.656 15.744 ;
  LAYER M1 ;
        RECT 30.624 16.176 30.656 16.92 ;
  LAYER M1 ;
        RECT 30.624 17.352 30.656 18.096 ;
  LAYER M1 ;
        RECT 30.624 18.528 30.656 19.272 ;
  LAYER M1 ;
        RECT 30.624 19.704 30.656 20.448 ;
  LAYER M1 ;
        RECT 30.624 20.88 30.656 21.624 ;
  LAYER M1 ;
        RECT 30.624 22.056 30.656 22.8 ;
  LAYER M1 ;
        RECT 30.624 23.232 30.656 23.976 ;
  LAYER M1 ;
        RECT 30.704 12.648 30.736 13.392 ;
  LAYER M1 ;
        RECT 30.704 13.488 30.736 13.728 ;
  LAYER M1 ;
        RECT 30.704 13.824 30.736 14.568 ;
  LAYER M1 ;
        RECT 30.704 14.664 30.736 14.904 ;
  LAYER M1 ;
        RECT 30.704 15 30.736 15.744 ;
  LAYER M1 ;
        RECT 30.704 15.84 30.736 16.08 ;
  LAYER M1 ;
        RECT 30.704 16.176 30.736 16.92 ;
  LAYER M1 ;
        RECT 30.704 17.016 30.736 17.256 ;
  LAYER M1 ;
        RECT 30.704 17.352 30.736 18.096 ;
  LAYER M1 ;
        RECT 30.704 18.192 30.736 18.432 ;
  LAYER M1 ;
        RECT 30.704 18.528 30.736 19.272 ;
  LAYER M1 ;
        RECT 30.704 19.368 30.736 19.608 ;
  LAYER M1 ;
        RECT 30.704 19.704 30.736 20.448 ;
  LAYER M1 ;
        RECT 30.704 20.544 30.736 20.784 ;
  LAYER M1 ;
        RECT 30.704 20.88 30.736 21.624 ;
  LAYER M1 ;
        RECT 30.704 21.72 30.736 21.96 ;
  LAYER M1 ;
        RECT 30.704 22.056 30.736 22.8 ;
  LAYER M1 ;
        RECT 30.704 22.896 30.736 23.136 ;
  LAYER M1 ;
        RECT 30.704 23.232 30.736 23.976 ;
  LAYER M1 ;
        RECT 30.704 24.072 30.736 24.312 ;
  LAYER M1 ;
        RECT 30.704 24.576 30.736 24.816 ;
  LAYER M1 ;
        RECT 30.784 12.648 30.816 13.392 ;
  LAYER M1 ;
        RECT 30.784 13.824 30.816 14.568 ;
  LAYER M1 ;
        RECT 30.784 15 30.816 15.744 ;
  LAYER M1 ;
        RECT 30.784 16.176 30.816 16.92 ;
  LAYER M1 ;
        RECT 30.784 17.352 30.816 18.096 ;
  LAYER M1 ;
        RECT 30.784 18.528 30.816 19.272 ;
  LAYER M1 ;
        RECT 30.784 19.704 30.816 20.448 ;
  LAYER M1 ;
        RECT 30.784 20.88 30.816 21.624 ;
  LAYER M1 ;
        RECT 30.784 22.056 30.816 22.8 ;
  LAYER M1 ;
        RECT 30.784 23.232 30.816 23.976 ;
  LAYER M1 ;
        RECT 30.864 12.648 30.896 13.392 ;
  LAYER M1 ;
        RECT 30.864 13.488 30.896 13.728 ;
  LAYER M1 ;
        RECT 30.864 13.824 30.896 14.568 ;
  LAYER M1 ;
        RECT 30.864 14.664 30.896 14.904 ;
  LAYER M1 ;
        RECT 30.864 15 30.896 15.744 ;
  LAYER M1 ;
        RECT 30.864 15.84 30.896 16.08 ;
  LAYER M1 ;
        RECT 30.864 16.176 30.896 16.92 ;
  LAYER M1 ;
        RECT 30.864 17.016 30.896 17.256 ;
  LAYER M1 ;
        RECT 30.864 17.352 30.896 18.096 ;
  LAYER M1 ;
        RECT 30.864 18.192 30.896 18.432 ;
  LAYER M1 ;
        RECT 30.864 18.528 30.896 19.272 ;
  LAYER M1 ;
        RECT 30.864 19.368 30.896 19.608 ;
  LAYER M1 ;
        RECT 30.864 19.704 30.896 20.448 ;
  LAYER M1 ;
        RECT 30.864 20.544 30.896 20.784 ;
  LAYER M1 ;
        RECT 30.864 20.88 30.896 21.624 ;
  LAYER M1 ;
        RECT 30.864 21.72 30.896 21.96 ;
  LAYER M1 ;
        RECT 30.864 22.056 30.896 22.8 ;
  LAYER M1 ;
        RECT 30.864 22.896 30.896 23.136 ;
  LAYER M1 ;
        RECT 30.864 23.232 30.896 23.976 ;
  LAYER M1 ;
        RECT 30.864 24.072 30.896 24.312 ;
  LAYER M1 ;
        RECT 30.864 24.576 30.896 24.816 ;
  LAYER M1 ;
        RECT 30.944 12.648 30.976 13.392 ;
  LAYER M1 ;
        RECT 30.944 13.824 30.976 14.568 ;
  LAYER M1 ;
        RECT 30.944 15 30.976 15.744 ;
  LAYER M1 ;
        RECT 30.944 16.176 30.976 16.92 ;
  LAYER M1 ;
        RECT 30.944 17.352 30.976 18.096 ;
  LAYER M1 ;
        RECT 30.944 18.528 30.976 19.272 ;
  LAYER M1 ;
        RECT 30.944 19.704 30.976 20.448 ;
  LAYER M1 ;
        RECT 30.944 20.88 30.976 21.624 ;
  LAYER M1 ;
        RECT 30.944 22.056 30.976 22.8 ;
  LAYER M1 ;
        RECT 30.944 23.232 30.976 23.976 ;
  LAYER M1 ;
        RECT 31.024 12.648 31.056 13.392 ;
  LAYER M1 ;
        RECT 31.024 13.488 31.056 13.728 ;
  LAYER M1 ;
        RECT 31.024 13.824 31.056 14.568 ;
  LAYER M1 ;
        RECT 31.024 14.664 31.056 14.904 ;
  LAYER M1 ;
        RECT 31.024 15 31.056 15.744 ;
  LAYER M1 ;
        RECT 31.024 15.84 31.056 16.08 ;
  LAYER M1 ;
        RECT 31.024 16.176 31.056 16.92 ;
  LAYER M1 ;
        RECT 31.024 17.016 31.056 17.256 ;
  LAYER M1 ;
        RECT 31.024 17.352 31.056 18.096 ;
  LAYER M1 ;
        RECT 31.024 18.192 31.056 18.432 ;
  LAYER M1 ;
        RECT 31.024 18.528 31.056 19.272 ;
  LAYER M1 ;
        RECT 31.024 19.368 31.056 19.608 ;
  LAYER M1 ;
        RECT 31.024 19.704 31.056 20.448 ;
  LAYER M1 ;
        RECT 31.024 20.544 31.056 20.784 ;
  LAYER M1 ;
        RECT 31.024 20.88 31.056 21.624 ;
  LAYER M1 ;
        RECT 31.024 21.72 31.056 21.96 ;
  LAYER M1 ;
        RECT 31.024 22.056 31.056 22.8 ;
  LAYER M1 ;
        RECT 31.024 22.896 31.056 23.136 ;
  LAYER M1 ;
        RECT 31.024 23.232 31.056 23.976 ;
  LAYER M1 ;
        RECT 31.024 24.072 31.056 24.312 ;
  LAYER M1 ;
        RECT 31.024 24.576 31.056 24.816 ;
  LAYER M1 ;
        RECT 31.104 12.648 31.136 13.392 ;
  LAYER M1 ;
        RECT 31.104 13.824 31.136 14.568 ;
  LAYER M1 ;
        RECT 31.104 15 31.136 15.744 ;
  LAYER M1 ;
        RECT 31.104 16.176 31.136 16.92 ;
  LAYER M1 ;
        RECT 31.104 17.352 31.136 18.096 ;
  LAYER M1 ;
        RECT 31.104 18.528 31.136 19.272 ;
  LAYER M1 ;
        RECT 31.104 19.704 31.136 20.448 ;
  LAYER M1 ;
        RECT 31.104 20.88 31.136 21.624 ;
  LAYER M1 ;
        RECT 31.104 22.056 31.136 22.8 ;
  LAYER M1 ;
        RECT 31.104 23.232 31.136 23.976 ;
  LAYER M1 ;
        RECT 31.184 12.648 31.216 13.392 ;
  LAYER M1 ;
        RECT 31.184 13.488 31.216 13.728 ;
  LAYER M1 ;
        RECT 31.184 13.824 31.216 14.568 ;
  LAYER M1 ;
        RECT 31.184 14.664 31.216 14.904 ;
  LAYER M1 ;
        RECT 31.184 15 31.216 15.744 ;
  LAYER M1 ;
        RECT 31.184 15.84 31.216 16.08 ;
  LAYER M1 ;
        RECT 31.184 16.176 31.216 16.92 ;
  LAYER M1 ;
        RECT 31.184 17.016 31.216 17.256 ;
  LAYER M1 ;
        RECT 31.184 17.352 31.216 18.096 ;
  LAYER M1 ;
        RECT 31.184 18.192 31.216 18.432 ;
  LAYER M1 ;
        RECT 31.184 18.528 31.216 19.272 ;
  LAYER M1 ;
        RECT 31.184 19.368 31.216 19.608 ;
  LAYER M1 ;
        RECT 31.184 19.704 31.216 20.448 ;
  LAYER M1 ;
        RECT 31.184 20.544 31.216 20.784 ;
  LAYER M1 ;
        RECT 31.184 20.88 31.216 21.624 ;
  LAYER M1 ;
        RECT 31.184 21.72 31.216 21.96 ;
  LAYER M1 ;
        RECT 31.184 22.056 31.216 22.8 ;
  LAYER M1 ;
        RECT 31.184 22.896 31.216 23.136 ;
  LAYER M1 ;
        RECT 31.184 23.232 31.216 23.976 ;
  LAYER M1 ;
        RECT 31.184 24.072 31.216 24.312 ;
  LAYER M1 ;
        RECT 31.184 24.576 31.216 24.816 ;
  LAYER M1 ;
        RECT 31.264 12.648 31.296 13.392 ;
  LAYER M1 ;
        RECT 31.264 13.824 31.296 14.568 ;
  LAYER M1 ;
        RECT 31.264 15 31.296 15.744 ;
  LAYER M1 ;
        RECT 31.264 16.176 31.296 16.92 ;
  LAYER M1 ;
        RECT 31.264 17.352 31.296 18.096 ;
  LAYER M1 ;
        RECT 31.264 18.528 31.296 19.272 ;
  LAYER M1 ;
        RECT 31.264 19.704 31.296 20.448 ;
  LAYER M1 ;
        RECT 31.264 20.88 31.296 21.624 ;
  LAYER M1 ;
        RECT 31.264 22.056 31.296 22.8 ;
  LAYER M1 ;
        RECT 31.264 23.232 31.296 23.976 ;
  LAYER M1 ;
        RECT 31.344 12.648 31.376 13.392 ;
  LAYER M1 ;
        RECT 31.344 13.488 31.376 13.728 ;
  LAYER M1 ;
        RECT 31.344 13.824 31.376 14.568 ;
  LAYER M1 ;
        RECT 31.344 14.664 31.376 14.904 ;
  LAYER M1 ;
        RECT 31.344 15 31.376 15.744 ;
  LAYER M1 ;
        RECT 31.344 15.84 31.376 16.08 ;
  LAYER M1 ;
        RECT 31.344 16.176 31.376 16.92 ;
  LAYER M1 ;
        RECT 31.344 17.016 31.376 17.256 ;
  LAYER M1 ;
        RECT 31.344 17.352 31.376 18.096 ;
  LAYER M1 ;
        RECT 31.344 18.192 31.376 18.432 ;
  LAYER M1 ;
        RECT 31.344 18.528 31.376 19.272 ;
  LAYER M1 ;
        RECT 31.344 19.368 31.376 19.608 ;
  LAYER M1 ;
        RECT 31.344 19.704 31.376 20.448 ;
  LAYER M1 ;
        RECT 31.344 20.544 31.376 20.784 ;
  LAYER M1 ;
        RECT 31.344 20.88 31.376 21.624 ;
  LAYER M1 ;
        RECT 31.344 21.72 31.376 21.96 ;
  LAYER M1 ;
        RECT 31.344 22.056 31.376 22.8 ;
  LAYER M1 ;
        RECT 31.344 22.896 31.376 23.136 ;
  LAYER M1 ;
        RECT 31.344 23.232 31.376 23.976 ;
  LAYER M1 ;
        RECT 31.344 24.072 31.376 24.312 ;
  LAYER M1 ;
        RECT 31.344 24.576 31.376 24.816 ;
  LAYER M1 ;
        RECT 31.424 12.648 31.456 13.392 ;
  LAYER M1 ;
        RECT 31.424 13.824 31.456 14.568 ;
  LAYER M1 ;
        RECT 31.424 15 31.456 15.744 ;
  LAYER M1 ;
        RECT 31.424 16.176 31.456 16.92 ;
  LAYER M1 ;
        RECT 31.424 17.352 31.456 18.096 ;
  LAYER M1 ;
        RECT 31.424 18.528 31.456 19.272 ;
  LAYER M1 ;
        RECT 31.424 19.704 31.456 20.448 ;
  LAYER M1 ;
        RECT 31.424 20.88 31.456 21.624 ;
  LAYER M1 ;
        RECT 31.424 22.056 31.456 22.8 ;
  LAYER M1 ;
        RECT 31.424 23.232 31.456 23.976 ;
  LAYER M1 ;
        RECT 31.504 12.648 31.536 13.392 ;
  LAYER M1 ;
        RECT 31.504 13.488 31.536 13.728 ;
  LAYER M1 ;
        RECT 31.504 13.824 31.536 14.568 ;
  LAYER M1 ;
        RECT 31.504 14.664 31.536 14.904 ;
  LAYER M1 ;
        RECT 31.504 15 31.536 15.744 ;
  LAYER M1 ;
        RECT 31.504 15.84 31.536 16.08 ;
  LAYER M1 ;
        RECT 31.504 16.176 31.536 16.92 ;
  LAYER M1 ;
        RECT 31.504 17.016 31.536 17.256 ;
  LAYER M1 ;
        RECT 31.504 17.352 31.536 18.096 ;
  LAYER M1 ;
        RECT 31.504 18.192 31.536 18.432 ;
  LAYER M1 ;
        RECT 31.504 18.528 31.536 19.272 ;
  LAYER M1 ;
        RECT 31.504 19.368 31.536 19.608 ;
  LAYER M1 ;
        RECT 31.504 19.704 31.536 20.448 ;
  LAYER M1 ;
        RECT 31.504 20.544 31.536 20.784 ;
  LAYER M1 ;
        RECT 31.504 20.88 31.536 21.624 ;
  LAYER M1 ;
        RECT 31.504 21.72 31.536 21.96 ;
  LAYER M1 ;
        RECT 31.504 22.056 31.536 22.8 ;
  LAYER M1 ;
        RECT 31.504 22.896 31.536 23.136 ;
  LAYER M1 ;
        RECT 31.504 23.232 31.536 23.976 ;
  LAYER M1 ;
        RECT 31.504 24.072 31.536 24.312 ;
  LAYER M1 ;
        RECT 31.504 24.576 31.536 24.816 ;
  LAYER M1 ;
        RECT 31.584 12.648 31.616 13.392 ;
  LAYER M1 ;
        RECT 31.584 13.824 31.616 14.568 ;
  LAYER M1 ;
        RECT 31.584 15 31.616 15.744 ;
  LAYER M1 ;
        RECT 31.584 16.176 31.616 16.92 ;
  LAYER M1 ;
        RECT 31.584 17.352 31.616 18.096 ;
  LAYER M1 ;
        RECT 31.584 18.528 31.616 19.272 ;
  LAYER M1 ;
        RECT 31.584 19.704 31.616 20.448 ;
  LAYER M1 ;
        RECT 31.584 20.88 31.616 21.624 ;
  LAYER M1 ;
        RECT 31.584 22.056 31.616 22.8 ;
  LAYER M1 ;
        RECT 31.584 23.232 31.616 23.976 ;
  LAYER M2 ;
        RECT 27.564 12.668 31.636 12.7 ;
  LAYER M2 ;
        RECT 27.644 12.752 31.556 12.784 ;
  LAYER M2 ;
        RECT 27.644 13.508 31.556 13.54 ;
  LAYER M2 ;
        RECT 27.564 13.844 31.636 13.876 ;
  LAYER M2 ;
        RECT 27.644 13.928 31.556 13.96 ;
  LAYER M2 ;
        RECT 27.644 14.684 31.556 14.716 ;
  LAYER M2 ;
        RECT 27.564 15.02 31.636 15.052 ;
  LAYER M2 ;
        RECT 27.644 15.104 31.556 15.136 ;
  LAYER M2 ;
        RECT 27.644 15.86 31.556 15.892 ;
  LAYER M2 ;
        RECT 27.564 16.196 31.636 16.228 ;
  LAYER M2 ;
        RECT 27.644 16.28 31.556 16.312 ;
  LAYER M2 ;
        RECT 27.644 17.036 31.556 17.068 ;
  LAYER M2 ;
        RECT 27.564 17.372 31.636 17.404 ;
  LAYER M2 ;
        RECT 27.644 17.456 31.556 17.488 ;
  LAYER M2 ;
        RECT 27.644 18.212 31.556 18.244 ;
  LAYER M2 ;
        RECT 27.564 18.548 31.636 18.58 ;
  LAYER M2 ;
        RECT 27.644 18.632 31.556 18.664 ;
  LAYER M2 ;
        RECT 27.644 19.388 31.556 19.42 ;
  LAYER M2 ;
        RECT 27.564 19.724 31.636 19.756 ;
  LAYER M2 ;
        RECT 27.644 19.808 31.556 19.84 ;
  LAYER M2 ;
        RECT 27.644 20.564 31.556 20.596 ;
  LAYER M2 ;
        RECT 27.564 20.9 31.636 20.932 ;
  LAYER M2 ;
        RECT 27.644 20.984 31.556 21.016 ;
  LAYER M2 ;
        RECT 27.644 21.74 31.556 21.772 ;
  LAYER M2 ;
        RECT 27.564 22.076 31.636 22.108 ;
  LAYER M2 ;
        RECT 27.644 22.16 31.556 22.192 ;
  LAYER M2 ;
        RECT 27.644 22.916 31.556 22.948 ;
  LAYER M2 ;
        RECT 27.564 23.252 31.636 23.284 ;
  LAYER M2 ;
        RECT 27.644 23.336 31.556 23.368 ;
  LAYER M2 ;
        RECT 27.644 24.092 31.556 24.124 ;
  LAYER M1 ;
        RECT 27.664 25.164 27.696 25.908 ;
  LAYER M1 ;
        RECT 27.664 26.004 27.696 26.244 ;
  LAYER M1 ;
        RECT 27.664 26.34 27.696 27.084 ;
  LAYER M1 ;
        RECT 27.664 27.18 27.696 27.42 ;
  LAYER M1 ;
        RECT 27.664 27.516 27.696 28.26 ;
  LAYER M1 ;
        RECT 27.664 28.356 27.696 28.596 ;
  LAYER M1 ;
        RECT 27.664 28.692 27.696 29.436 ;
  LAYER M1 ;
        RECT 27.664 29.532 27.696 29.772 ;
  LAYER M1 ;
        RECT 27.664 29.868 27.696 30.612 ;
  LAYER M1 ;
        RECT 27.664 30.708 27.696 30.948 ;
  LAYER M1 ;
        RECT 27.664 31.044 27.696 31.788 ;
  LAYER M1 ;
        RECT 27.664 31.884 27.696 32.124 ;
  LAYER M1 ;
        RECT 27.664 32.22 27.696 32.964 ;
  LAYER M1 ;
        RECT 27.664 33.06 27.696 33.3 ;
  LAYER M1 ;
        RECT 27.664 33.396 27.696 34.14 ;
  LAYER M1 ;
        RECT 27.664 34.236 27.696 34.476 ;
  LAYER M1 ;
        RECT 27.664 34.572 27.696 35.316 ;
  LAYER M1 ;
        RECT 27.664 35.412 27.696 35.652 ;
  LAYER M1 ;
        RECT 27.664 35.748 27.696 36.492 ;
  LAYER M1 ;
        RECT 27.664 36.588 27.696 36.828 ;
  LAYER M1 ;
        RECT 27.664 37.092 27.696 37.332 ;
  LAYER M1 ;
        RECT 27.584 25.164 27.616 25.908 ;
  LAYER M1 ;
        RECT 27.584 26.34 27.616 27.084 ;
  LAYER M1 ;
        RECT 27.584 27.516 27.616 28.26 ;
  LAYER M1 ;
        RECT 27.584 28.692 27.616 29.436 ;
  LAYER M1 ;
        RECT 27.584 29.868 27.616 30.612 ;
  LAYER M1 ;
        RECT 27.584 31.044 27.616 31.788 ;
  LAYER M1 ;
        RECT 27.584 32.22 27.616 32.964 ;
  LAYER M1 ;
        RECT 27.584 33.396 27.616 34.14 ;
  LAYER M1 ;
        RECT 27.584 34.572 27.616 35.316 ;
  LAYER M1 ;
        RECT 27.584 35.748 27.616 36.492 ;
  LAYER M1 ;
        RECT 27.744 25.164 27.776 25.908 ;
  LAYER M1 ;
        RECT 27.744 26.34 27.776 27.084 ;
  LAYER M1 ;
        RECT 27.744 27.516 27.776 28.26 ;
  LAYER M1 ;
        RECT 27.744 28.692 27.776 29.436 ;
  LAYER M1 ;
        RECT 27.744 29.868 27.776 30.612 ;
  LAYER M1 ;
        RECT 27.744 31.044 27.776 31.788 ;
  LAYER M1 ;
        RECT 27.744 32.22 27.776 32.964 ;
  LAYER M1 ;
        RECT 27.744 33.396 27.776 34.14 ;
  LAYER M1 ;
        RECT 27.744 34.572 27.776 35.316 ;
  LAYER M1 ;
        RECT 27.744 35.748 27.776 36.492 ;
  LAYER M1 ;
        RECT 27.824 25.164 27.856 25.908 ;
  LAYER M1 ;
        RECT 27.824 26.004 27.856 26.244 ;
  LAYER M1 ;
        RECT 27.824 26.34 27.856 27.084 ;
  LAYER M1 ;
        RECT 27.824 27.18 27.856 27.42 ;
  LAYER M1 ;
        RECT 27.824 27.516 27.856 28.26 ;
  LAYER M1 ;
        RECT 27.824 28.356 27.856 28.596 ;
  LAYER M1 ;
        RECT 27.824 28.692 27.856 29.436 ;
  LAYER M1 ;
        RECT 27.824 29.532 27.856 29.772 ;
  LAYER M1 ;
        RECT 27.824 29.868 27.856 30.612 ;
  LAYER M1 ;
        RECT 27.824 30.708 27.856 30.948 ;
  LAYER M1 ;
        RECT 27.824 31.044 27.856 31.788 ;
  LAYER M1 ;
        RECT 27.824 31.884 27.856 32.124 ;
  LAYER M1 ;
        RECT 27.824 32.22 27.856 32.964 ;
  LAYER M1 ;
        RECT 27.824 33.06 27.856 33.3 ;
  LAYER M1 ;
        RECT 27.824 33.396 27.856 34.14 ;
  LAYER M1 ;
        RECT 27.824 34.236 27.856 34.476 ;
  LAYER M1 ;
        RECT 27.824 34.572 27.856 35.316 ;
  LAYER M1 ;
        RECT 27.824 35.412 27.856 35.652 ;
  LAYER M1 ;
        RECT 27.824 35.748 27.856 36.492 ;
  LAYER M1 ;
        RECT 27.824 36.588 27.856 36.828 ;
  LAYER M1 ;
        RECT 27.824 37.092 27.856 37.332 ;
  LAYER M1 ;
        RECT 27.904 25.164 27.936 25.908 ;
  LAYER M1 ;
        RECT 27.904 26.34 27.936 27.084 ;
  LAYER M1 ;
        RECT 27.904 27.516 27.936 28.26 ;
  LAYER M1 ;
        RECT 27.904 28.692 27.936 29.436 ;
  LAYER M1 ;
        RECT 27.904 29.868 27.936 30.612 ;
  LAYER M1 ;
        RECT 27.904 31.044 27.936 31.788 ;
  LAYER M1 ;
        RECT 27.904 32.22 27.936 32.964 ;
  LAYER M1 ;
        RECT 27.904 33.396 27.936 34.14 ;
  LAYER M1 ;
        RECT 27.904 34.572 27.936 35.316 ;
  LAYER M1 ;
        RECT 27.904 35.748 27.936 36.492 ;
  LAYER M1 ;
        RECT 27.984 25.164 28.016 25.908 ;
  LAYER M1 ;
        RECT 27.984 26.004 28.016 26.244 ;
  LAYER M1 ;
        RECT 27.984 26.34 28.016 27.084 ;
  LAYER M1 ;
        RECT 27.984 27.18 28.016 27.42 ;
  LAYER M1 ;
        RECT 27.984 27.516 28.016 28.26 ;
  LAYER M1 ;
        RECT 27.984 28.356 28.016 28.596 ;
  LAYER M1 ;
        RECT 27.984 28.692 28.016 29.436 ;
  LAYER M1 ;
        RECT 27.984 29.532 28.016 29.772 ;
  LAYER M1 ;
        RECT 27.984 29.868 28.016 30.612 ;
  LAYER M1 ;
        RECT 27.984 30.708 28.016 30.948 ;
  LAYER M1 ;
        RECT 27.984 31.044 28.016 31.788 ;
  LAYER M1 ;
        RECT 27.984 31.884 28.016 32.124 ;
  LAYER M1 ;
        RECT 27.984 32.22 28.016 32.964 ;
  LAYER M1 ;
        RECT 27.984 33.06 28.016 33.3 ;
  LAYER M1 ;
        RECT 27.984 33.396 28.016 34.14 ;
  LAYER M1 ;
        RECT 27.984 34.236 28.016 34.476 ;
  LAYER M1 ;
        RECT 27.984 34.572 28.016 35.316 ;
  LAYER M1 ;
        RECT 27.984 35.412 28.016 35.652 ;
  LAYER M1 ;
        RECT 27.984 35.748 28.016 36.492 ;
  LAYER M1 ;
        RECT 27.984 36.588 28.016 36.828 ;
  LAYER M1 ;
        RECT 27.984 37.092 28.016 37.332 ;
  LAYER M1 ;
        RECT 28.064 25.164 28.096 25.908 ;
  LAYER M1 ;
        RECT 28.064 26.34 28.096 27.084 ;
  LAYER M1 ;
        RECT 28.064 27.516 28.096 28.26 ;
  LAYER M1 ;
        RECT 28.064 28.692 28.096 29.436 ;
  LAYER M1 ;
        RECT 28.064 29.868 28.096 30.612 ;
  LAYER M1 ;
        RECT 28.064 31.044 28.096 31.788 ;
  LAYER M1 ;
        RECT 28.064 32.22 28.096 32.964 ;
  LAYER M1 ;
        RECT 28.064 33.396 28.096 34.14 ;
  LAYER M1 ;
        RECT 28.064 34.572 28.096 35.316 ;
  LAYER M1 ;
        RECT 28.064 35.748 28.096 36.492 ;
  LAYER M1 ;
        RECT 28.144 25.164 28.176 25.908 ;
  LAYER M1 ;
        RECT 28.144 26.004 28.176 26.244 ;
  LAYER M1 ;
        RECT 28.144 26.34 28.176 27.084 ;
  LAYER M1 ;
        RECT 28.144 27.18 28.176 27.42 ;
  LAYER M1 ;
        RECT 28.144 27.516 28.176 28.26 ;
  LAYER M1 ;
        RECT 28.144 28.356 28.176 28.596 ;
  LAYER M1 ;
        RECT 28.144 28.692 28.176 29.436 ;
  LAYER M1 ;
        RECT 28.144 29.532 28.176 29.772 ;
  LAYER M1 ;
        RECT 28.144 29.868 28.176 30.612 ;
  LAYER M1 ;
        RECT 28.144 30.708 28.176 30.948 ;
  LAYER M1 ;
        RECT 28.144 31.044 28.176 31.788 ;
  LAYER M1 ;
        RECT 28.144 31.884 28.176 32.124 ;
  LAYER M1 ;
        RECT 28.144 32.22 28.176 32.964 ;
  LAYER M1 ;
        RECT 28.144 33.06 28.176 33.3 ;
  LAYER M1 ;
        RECT 28.144 33.396 28.176 34.14 ;
  LAYER M1 ;
        RECT 28.144 34.236 28.176 34.476 ;
  LAYER M1 ;
        RECT 28.144 34.572 28.176 35.316 ;
  LAYER M1 ;
        RECT 28.144 35.412 28.176 35.652 ;
  LAYER M1 ;
        RECT 28.144 35.748 28.176 36.492 ;
  LAYER M1 ;
        RECT 28.144 36.588 28.176 36.828 ;
  LAYER M1 ;
        RECT 28.144 37.092 28.176 37.332 ;
  LAYER M1 ;
        RECT 28.224 25.164 28.256 25.908 ;
  LAYER M1 ;
        RECT 28.224 26.34 28.256 27.084 ;
  LAYER M1 ;
        RECT 28.224 27.516 28.256 28.26 ;
  LAYER M1 ;
        RECT 28.224 28.692 28.256 29.436 ;
  LAYER M1 ;
        RECT 28.224 29.868 28.256 30.612 ;
  LAYER M1 ;
        RECT 28.224 31.044 28.256 31.788 ;
  LAYER M1 ;
        RECT 28.224 32.22 28.256 32.964 ;
  LAYER M1 ;
        RECT 28.224 33.396 28.256 34.14 ;
  LAYER M1 ;
        RECT 28.224 34.572 28.256 35.316 ;
  LAYER M1 ;
        RECT 28.224 35.748 28.256 36.492 ;
  LAYER M1 ;
        RECT 28.304 25.164 28.336 25.908 ;
  LAYER M1 ;
        RECT 28.304 26.004 28.336 26.244 ;
  LAYER M1 ;
        RECT 28.304 26.34 28.336 27.084 ;
  LAYER M1 ;
        RECT 28.304 27.18 28.336 27.42 ;
  LAYER M1 ;
        RECT 28.304 27.516 28.336 28.26 ;
  LAYER M1 ;
        RECT 28.304 28.356 28.336 28.596 ;
  LAYER M1 ;
        RECT 28.304 28.692 28.336 29.436 ;
  LAYER M1 ;
        RECT 28.304 29.532 28.336 29.772 ;
  LAYER M1 ;
        RECT 28.304 29.868 28.336 30.612 ;
  LAYER M1 ;
        RECT 28.304 30.708 28.336 30.948 ;
  LAYER M1 ;
        RECT 28.304 31.044 28.336 31.788 ;
  LAYER M1 ;
        RECT 28.304 31.884 28.336 32.124 ;
  LAYER M1 ;
        RECT 28.304 32.22 28.336 32.964 ;
  LAYER M1 ;
        RECT 28.304 33.06 28.336 33.3 ;
  LAYER M1 ;
        RECT 28.304 33.396 28.336 34.14 ;
  LAYER M1 ;
        RECT 28.304 34.236 28.336 34.476 ;
  LAYER M1 ;
        RECT 28.304 34.572 28.336 35.316 ;
  LAYER M1 ;
        RECT 28.304 35.412 28.336 35.652 ;
  LAYER M1 ;
        RECT 28.304 35.748 28.336 36.492 ;
  LAYER M1 ;
        RECT 28.304 36.588 28.336 36.828 ;
  LAYER M1 ;
        RECT 28.304 37.092 28.336 37.332 ;
  LAYER M1 ;
        RECT 28.384 25.164 28.416 25.908 ;
  LAYER M1 ;
        RECT 28.384 26.34 28.416 27.084 ;
  LAYER M1 ;
        RECT 28.384 27.516 28.416 28.26 ;
  LAYER M1 ;
        RECT 28.384 28.692 28.416 29.436 ;
  LAYER M1 ;
        RECT 28.384 29.868 28.416 30.612 ;
  LAYER M1 ;
        RECT 28.384 31.044 28.416 31.788 ;
  LAYER M1 ;
        RECT 28.384 32.22 28.416 32.964 ;
  LAYER M1 ;
        RECT 28.384 33.396 28.416 34.14 ;
  LAYER M1 ;
        RECT 28.384 34.572 28.416 35.316 ;
  LAYER M1 ;
        RECT 28.384 35.748 28.416 36.492 ;
  LAYER M1 ;
        RECT 28.464 25.164 28.496 25.908 ;
  LAYER M1 ;
        RECT 28.464 26.004 28.496 26.244 ;
  LAYER M1 ;
        RECT 28.464 26.34 28.496 27.084 ;
  LAYER M1 ;
        RECT 28.464 27.18 28.496 27.42 ;
  LAYER M1 ;
        RECT 28.464 27.516 28.496 28.26 ;
  LAYER M1 ;
        RECT 28.464 28.356 28.496 28.596 ;
  LAYER M1 ;
        RECT 28.464 28.692 28.496 29.436 ;
  LAYER M1 ;
        RECT 28.464 29.532 28.496 29.772 ;
  LAYER M1 ;
        RECT 28.464 29.868 28.496 30.612 ;
  LAYER M1 ;
        RECT 28.464 30.708 28.496 30.948 ;
  LAYER M1 ;
        RECT 28.464 31.044 28.496 31.788 ;
  LAYER M1 ;
        RECT 28.464 31.884 28.496 32.124 ;
  LAYER M1 ;
        RECT 28.464 32.22 28.496 32.964 ;
  LAYER M1 ;
        RECT 28.464 33.06 28.496 33.3 ;
  LAYER M1 ;
        RECT 28.464 33.396 28.496 34.14 ;
  LAYER M1 ;
        RECT 28.464 34.236 28.496 34.476 ;
  LAYER M1 ;
        RECT 28.464 34.572 28.496 35.316 ;
  LAYER M1 ;
        RECT 28.464 35.412 28.496 35.652 ;
  LAYER M1 ;
        RECT 28.464 35.748 28.496 36.492 ;
  LAYER M1 ;
        RECT 28.464 36.588 28.496 36.828 ;
  LAYER M1 ;
        RECT 28.464 37.092 28.496 37.332 ;
  LAYER M1 ;
        RECT 28.544 25.164 28.576 25.908 ;
  LAYER M1 ;
        RECT 28.544 26.34 28.576 27.084 ;
  LAYER M1 ;
        RECT 28.544 27.516 28.576 28.26 ;
  LAYER M1 ;
        RECT 28.544 28.692 28.576 29.436 ;
  LAYER M1 ;
        RECT 28.544 29.868 28.576 30.612 ;
  LAYER M1 ;
        RECT 28.544 31.044 28.576 31.788 ;
  LAYER M1 ;
        RECT 28.544 32.22 28.576 32.964 ;
  LAYER M1 ;
        RECT 28.544 33.396 28.576 34.14 ;
  LAYER M1 ;
        RECT 28.544 34.572 28.576 35.316 ;
  LAYER M1 ;
        RECT 28.544 35.748 28.576 36.492 ;
  LAYER M1 ;
        RECT 28.624 25.164 28.656 25.908 ;
  LAYER M1 ;
        RECT 28.624 26.004 28.656 26.244 ;
  LAYER M1 ;
        RECT 28.624 26.34 28.656 27.084 ;
  LAYER M1 ;
        RECT 28.624 27.18 28.656 27.42 ;
  LAYER M1 ;
        RECT 28.624 27.516 28.656 28.26 ;
  LAYER M1 ;
        RECT 28.624 28.356 28.656 28.596 ;
  LAYER M1 ;
        RECT 28.624 28.692 28.656 29.436 ;
  LAYER M1 ;
        RECT 28.624 29.532 28.656 29.772 ;
  LAYER M1 ;
        RECT 28.624 29.868 28.656 30.612 ;
  LAYER M1 ;
        RECT 28.624 30.708 28.656 30.948 ;
  LAYER M1 ;
        RECT 28.624 31.044 28.656 31.788 ;
  LAYER M1 ;
        RECT 28.624 31.884 28.656 32.124 ;
  LAYER M1 ;
        RECT 28.624 32.22 28.656 32.964 ;
  LAYER M1 ;
        RECT 28.624 33.06 28.656 33.3 ;
  LAYER M1 ;
        RECT 28.624 33.396 28.656 34.14 ;
  LAYER M1 ;
        RECT 28.624 34.236 28.656 34.476 ;
  LAYER M1 ;
        RECT 28.624 34.572 28.656 35.316 ;
  LAYER M1 ;
        RECT 28.624 35.412 28.656 35.652 ;
  LAYER M1 ;
        RECT 28.624 35.748 28.656 36.492 ;
  LAYER M1 ;
        RECT 28.624 36.588 28.656 36.828 ;
  LAYER M1 ;
        RECT 28.624 37.092 28.656 37.332 ;
  LAYER M1 ;
        RECT 28.704 25.164 28.736 25.908 ;
  LAYER M1 ;
        RECT 28.704 26.34 28.736 27.084 ;
  LAYER M1 ;
        RECT 28.704 27.516 28.736 28.26 ;
  LAYER M1 ;
        RECT 28.704 28.692 28.736 29.436 ;
  LAYER M1 ;
        RECT 28.704 29.868 28.736 30.612 ;
  LAYER M1 ;
        RECT 28.704 31.044 28.736 31.788 ;
  LAYER M1 ;
        RECT 28.704 32.22 28.736 32.964 ;
  LAYER M1 ;
        RECT 28.704 33.396 28.736 34.14 ;
  LAYER M1 ;
        RECT 28.704 34.572 28.736 35.316 ;
  LAYER M1 ;
        RECT 28.704 35.748 28.736 36.492 ;
  LAYER M1 ;
        RECT 28.784 25.164 28.816 25.908 ;
  LAYER M1 ;
        RECT 28.784 26.004 28.816 26.244 ;
  LAYER M1 ;
        RECT 28.784 26.34 28.816 27.084 ;
  LAYER M1 ;
        RECT 28.784 27.18 28.816 27.42 ;
  LAYER M1 ;
        RECT 28.784 27.516 28.816 28.26 ;
  LAYER M1 ;
        RECT 28.784 28.356 28.816 28.596 ;
  LAYER M1 ;
        RECT 28.784 28.692 28.816 29.436 ;
  LAYER M1 ;
        RECT 28.784 29.532 28.816 29.772 ;
  LAYER M1 ;
        RECT 28.784 29.868 28.816 30.612 ;
  LAYER M1 ;
        RECT 28.784 30.708 28.816 30.948 ;
  LAYER M1 ;
        RECT 28.784 31.044 28.816 31.788 ;
  LAYER M1 ;
        RECT 28.784 31.884 28.816 32.124 ;
  LAYER M1 ;
        RECT 28.784 32.22 28.816 32.964 ;
  LAYER M1 ;
        RECT 28.784 33.06 28.816 33.3 ;
  LAYER M1 ;
        RECT 28.784 33.396 28.816 34.14 ;
  LAYER M1 ;
        RECT 28.784 34.236 28.816 34.476 ;
  LAYER M1 ;
        RECT 28.784 34.572 28.816 35.316 ;
  LAYER M1 ;
        RECT 28.784 35.412 28.816 35.652 ;
  LAYER M1 ;
        RECT 28.784 35.748 28.816 36.492 ;
  LAYER M1 ;
        RECT 28.784 36.588 28.816 36.828 ;
  LAYER M1 ;
        RECT 28.784 37.092 28.816 37.332 ;
  LAYER M1 ;
        RECT 28.864 25.164 28.896 25.908 ;
  LAYER M1 ;
        RECT 28.864 26.34 28.896 27.084 ;
  LAYER M1 ;
        RECT 28.864 27.516 28.896 28.26 ;
  LAYER M1 ;
        RECT 28.864 28.692 28.896 29.436 ;
  LAYER M1 ;
        RECT 28.864 29.868 28.896 30.612 ;
  LAYER M1 ;
        RECT 28.864 31.044 28.896 31.788 ;
  LAYER M1 ;
        RECT 28.864 32.22 28.896 32.964 ;
  LAYER M1 ;
        RECT 28.864 33.396 28.896 34.14 ;
  LAYER M1 ;
        RECT 28.864 34.572 28.896 35.316 ;
  LAYER M1 ;
        RECT 28.864 35.748 28.896 36.492 ;
  LAYER M1 ;
        RECT 28.944 25.164 28.976 25.908 ;
  LAYER M1 ;
        RECT 28.944 26.004 28.976 26.244 ;
  LAYER M1 ;
        RECT 28.944 26.34 28.976 27.084 ;
  LAYER M1 ;
        RECT 28.944 27.18 28.976 27.42 ;
  LAYER M1 ;
        RECT 28.944 27.516 28.976 28.26 ;
  LAYER M1 ;
        RECT 28.944 28.356 28.976 28.596 ;
  LAYER M1 ;
        RECT 28.944 28.692 28.976 29.436 ;
  LAYER M1 ;
        RECT 28.944 29.532 28.976 29.772 ;
  LAYER M1 ;
        RECT 28.944 29.868 28.976 30.612 ;
  LAYER M1 ;
        RECT 28.944 30.708 28.976 30.948 ;
  LAYER M1 ;
        RECT 28.944 31.044 28.976 31.788 ;
  LAYER M1 ;
        RECT 28.944 31.884 28.976 32.124 ;
  LAYER M1 ;
        RECT 28.944 32.22 28.976 32.964 ;
  LAYER M1 ;
        RECT 28.944 33.06 28.976 33.3 ;
  LAYER M1 ;
        RECT 28.944 33.396 28.976 34.14 ;
  LAYER M1 ;
        RECT 28.944 34.236 28.976 34.476 ;
  LAYER M1 ;
        RECT 28.944 34.572 28.976 35.316 ;
  LAYER M1 ;
        RECT 28.944 35.412 28.976 35.652 ;
  LAYER M1 ;
        RECT 28.944 35.748 28.976 36.492 ;
  LAYER M1 ;
        RECT 28.944 36.588 28.976 36.828 ;
  LAYER M1 ;
        RECT 28.944 37.092 28.976 37.332 ;
  LAYER M1 ;
        RECT 29.024 25.164 29.056 25.908 ;
  LAYER M1 ;
        RECT 29.024 26.34 29.056 27.084 ;
  LAYER M1 ;
        RECT 29.024 27.516 29.056 28.26 ;
  LAYER M1 ;
        RECT 29.024 28.692 29.056 29.436 ;
  LAYER M1 ;
        RECT 29.024 29.868 29.056 30.612 ;
  LAYER M1 ;
        RECT 29.024 31.044 29.056 31.788 ;
  LAYER M1 ;
        RECT 29.024 32.22 29.056 32.964 ;
  LAYER M1 ;
        RECT 29.024 33.396 29.056 34.14 ;
  LAYER M1 ;
        RECT 29.024 34.572 29.056 35.316 ;
  LAYER M1 ;
        RECT 29.024 35.748 29.056 36.492 ;
  LAYER M1 ;
        RECT 29.104 25.164 29.136 25.908 ;
  LAYER M1 ;
        RECT 29.104 26.004 29.136 26.244 ;
  LAYER M1 ;
        RECT 29.104 26.34 29.136 27.084 ;
  LAYER M1 ;
        RECT 29.104 27.18 29.136 27.42 ;
  LAYER M1 ;
        RECT 29.104 27.516 29.136 28.26 ;
  LAYER M1 ;
        RECT 29.104 28.356 29.136 28.596 ;
  LAYER M1 ;
        RECT 29.104 28.692 29.136 29.436 ;
  LAYER M1 ;
        RECT 29.104 29.532 29.136 29.772 ;
  LAYER M1 ;
        RECT 29.104 29.868 29.136 30.612 ;
  LAYER M1 ;
        RECT 29.104 30.708 29.136 30.948 ;
  LAYER M1 ;
        RECT 29.104 31.044 29.136 31.788 ;
  LAYER M1 ;
        RECT 29.104 31.884 29.136 32.124 ;
  LAYER M1 ;
        RECT 29.104 32.22 29.136 32.964 ;
  LAYER M1 ;
        RECT 29.104 33.06 29.136 33.3 ;
  LAYER M1 ;
        RECT 29.104 33.396 29.136 34.14 ;
  LAYER M1 ;
        RECT 29.104 34.236 29.136 34.476 ;
  LAYER M1 ;
        RECT 29.104 34.572 29.136 35.316 ;
  LAYER M1 ;
        RECT 29.104 35.412 29.136 35.652 ;
  LAYER M1 ;
        RECT 29.104 35.748 29.136 36.492 ;
  LAYER M1 ;
        RECT 29.104 36.588 29.136 36.828 ;
  LAYER M1 ;
        RECT 29.104 37.092 29.136 37.332 ;
  LAYER M1 ;
        RECT 29.184 25.164 29.216 25.908 ;
  LAYER M1 ;
        RECT 29.184 26.34 29.216 27.084 ;
  LAYER M1 ;
        RECT 29.184 27.516 29.216 28.26 ;
  LAYER M1 ;
        RECT 29.184 28.692 29.216 29.436 ;
  LAYER M1 ;
        RECT 29.184 29.868 29.216 30.612 ;
  LAYER M1 ;
        RECT 29.184 31.044 29.216 31.788 ;
  LAYER M1 ;
        RECT 29.184 32.22 29.216 32.964 ;
  LAYER M1 ;
        RECT 29.184 33.396 29.216 34.14 ;
  LAYER M1 ;
        RECT 29.184 34.572 29.216 35.316 ;
  LAYER M1 ;
        RECT 29.184 35.748 29.216 36.492 ;
  LAYER M1 ;
        RECT 29.264 25.164 29.296 25.908 ;
  LAYER M1 ;
        RECT 29.264 26.004 29.296 26.244 ;
  LAYER M1 ;
        RECT 29.264 26.34 29.296 27.084 ;
  LAYER M1 ;
        RECT 29.264 27.18 29.296 27.42 ;
  LAYER M1 ;
        RECT 29.264 27.516 29.296 28.26 ;
  LAYER M1 ;
        RECT 29.264 28.356 29.296 28.596 ;
  LAYER M1 ;
        RECT 29.264 28.692 29.296 29.436 ;
  LAYER M1 ;
        RECT 29.264 29.532 29.296 29.772 ;
  LAYER M1 ;
        RECT 29.264 29.868 29.296 30.612 ;
  LAYER M1 ;
        RECT 29.264 30.708 29.296 30.948 ;
  LAYER M1 ;
        RECT 29.264 31.044 29.296 31.788 ;
  LAYER M1 ;
        RECT 29.264 31.884 29.296 32.124 ;
  LAYER M1 ;
        RECT 29.264 32.22 29.296 32.964 ;
  LAYER M1 ;
        RECT 29.264 33.06 29.296 33.3 ;
  LAYER M1 ;
        RECT 29.264 33.396 29.296 34.14 ;
  LAYER M1 ;
        RECT 29.264 34.236 29.296 34.476 ;
  LAYER M1 ;
        RECT 29.264 34.572 29.296 35.316 ;
  LAYER M1 ;
        RECT 29.264 35.412 29.296 35.652 ;
  LAYER M1 ;
        RECT 29.264 35.748 29.296 36.492 ;
  LAYER M1 ;
        RECT 29.264 36.588 29.296 36.828 ;
  LAYER M1 ;
        RECT 29.264 37.092 29.296 37.332 ;
  LAYER M1 ;
        RECT 29.344 25.164 29.376 25.908 ;
  LAYER M1 ;
        RECT 29.344 26.34 29.376 27.084 ;
  LAYER M1 ;
        RECT 29.344 27.516 29.376 28.26 ;
  LAYER M1 ;
        RECT 29.344 28.692 29.376 29.436 ;
  LAYER M1 ;
        RECT 29.344 29.868 29.376 30.612 ;
  LAYER M1 ;
        RECT 29.344 31.044 29.376 31.788 ;
  LAYER M1 ;
        RECT 29.344 32.22 29.376 32.964 ;
  LAYER M1 ;
        RECT 29.344 33.396 29.376 34.14 ;
  LAYER M1 ;
        RECT 29.344 34.572 29.376 35.316 ;
  LAYER M1 ;
        RECT 29.344 35.748 29.376 36.492 ;
  LAYER M1 ;
        RECT 29.424 25.164 29.456 25.908 ;
  LAYER M1 ;
        RECT 29.424 26.004 29.456 26.244 ;
  LAYER M1 ;
        RECT 29.424 26.34 29.456 27.084 ;
  LAYER M1 ;
        RECT 29.424 27.18 29.456 27.42 ;
  LAYER M1 ;
        RECT 29.424 27.516 29.456 28.26 ;
  LAYER M1 ;
        RECT 29.424 28.356 29.456 28.596 ;
  LAYER M1 ;
        RECT 29.424 28.692 29.456 29.436 ;
  LAYER M1 ;
        RECT 29.424 29.532 29.456 29.772 ;
  LAYER M1 ;
        RECT 29.424 29.868 29.456 30.612 ;
  LAYER M1 ;
        RECT 29.424 30.708 29.456 30.948 ;
  LAYER M1 ;
        RECT 29.424 31.044 29.456 31.788 ;
  LAYER M1 ;
        RECT 29.424 31.884 29.456 32.124 ;
  LAYER M1 ;
        RECT 29.424 32.22 29.456 32.964 ;
  LAYER M1 ;
        RECT 29.424 33.06 29.456 33.3 ;
  LAYER M1 ;
        RECT 29.424 33.396 29.456 34.14 ;
  LAYER M1 ;
        RECT 29.424 34.236 29.456 34.476 ;
  LAYER M1 ;
        RECT 29.424 34.572 29.456 35.316 ;
  LAYER M1 ;
        RECT 29.424 35.412 29.456 35.652 ;
  LAYER M1 ;
        RECT 29.424 35.748 29.456 36.492 ;
  LAYER M1 ;
        RECT 29.424 36.588 29.456 36.828 ;
  LAYER M1 ;
        RECT 29.424 37.092 29.456 37.332 ;
  LAYER M1 ;
        RECT 29.504 25.164 29.536 25.908 ;
  LAYER M1 ;
        RECT 29.504 26.34 29.536 27.084 ;
  LAYER M1 ;
        RECT 29.504 27.516 29.536 28.26 ;
  LAYER M1 ;
        RECT 29.504 28.692 29.536 29.436 ;
  LAYER M1 ;
        RECT 29.504 29.868 29.536 30.612 ;
  LAYER M1 ;
        RECT 29.504 31.044 29.536 31.788 ;
  LAYER M1 ;
        RECT 29.504 32.22 29.536 32.964 ;
  LAYER M1 ;
        RECT 29.504 33.396 29.536 34.14 ;
  LAYER M1 ;
        RECT 29.504 34.572 29.536 35.316 ;
  LAYER M1 ;
        RECT 29.504 35.748 29.536 36.492 ;
  LAYER M1 ;
        RECT 29.584 25.164 29.616 25.908 ;
  LAYER M1 ;
        RECT 29.584 26.004 29.616 26.244 ;
  LAYER M1 ;
        RECT 29.584 26.34 29.616 27.084 ;
  LAYER M1 ;
        RECT 29.584 27.18 29.616 27.42 ;
  LAYER M1 ;
        RECT 29.584 27.516 29.616 28.26 ;
  LAYER M1 ;
        RECT 29.584 28.356 29.616 28.596 ;
  LAYER M1 ;
        RECT 29.584 28.692 29.616 29.436 ;
  LAYER M1 ;
        RECT 29.584 29.532 29.616 29.772 ;
  LAYER M1 ;
        RECT 29.584 29.868 29.616 30.612 ;
  LAYER M1 ;
        RECT 29.584 30.708 29.616 30.948 ;
  LAYER M1 ;
        RECT 29.584 31.044 29.616 31.788 ;
  LAYER M1 ;
        RECT 29.584 31.884 29.616 32.124 ;
  LAYER M1 ;
        RECT 29.584 32.22 29.616 32.964 ;
  LAYER M1 ;
        RECT 29.584 33.06 29.616 33.3 ;
  LAYER M1 ;
        RECT 29.584 33.396 29.616 34.14 ;
  LAYER M1 ;
        RECT 29.584 34.236 29.616 34.476 ;
  LAYER M1 ;
        RECT 29.584 34.572 29.616 35.316 ;
  LAYER M1 ;
        RECT 29.584 35.412 29.616 35.652 ;
  LAYER M1 ;
        RECT 29.584 35.748 29.616 36.492 ;
  LAYER M1 ;
        RECT 29.584 36.588 29.616 36.828 ;
  LAYER M1 ;
        RECT 29.584 37.092 29.616 37.332 ;
  LAYER M1 ;
        RECT 29.664 25.164 29.696 25.908 ;
  LAYER M1 ;
        RECT 29.664 26.34 29.696 27.084 ;
  LAYER M1 ;
        RECT 29.664 27.516 29.696 28.26 ;
  LAYER M1 ;
        RECT 29.664 28.692 29.696 29.436 ;
  LAYER M1 ;
        RECT 29.664 29.868 29.696 30.612 ;
  LAYER M1 ;
        RECT 29.664 31.044 29.696 31.788 ;
  LAYER M1 ;
        RECT 29.664 32.22 29.696 32.964 ;
  LAYER M1 ;
        RECT 29.664 33.396 29.696 34.14 ;
  LAYER M1 ;
        RECT 29.664 34.572 29.696 35.316 ;
  LAYER M1 ;
        RECT 29.664 35.748 29.696 36.492 ;
  LAYER M1 ;
        RECT 29.744 25.164 29.776 25.908 ;
  LAYER M1 ;
        RECT 29.744 26.004 29.776 26.244 ;
  LAYER M1 ;
        RECT 29.744 26.34 29.776 27.084 ;
  LAYER M1 ;
        RECT 29.744 27.18 29.776 27.42 ;
  LAYER M1 ;
        RECT 29.744 27.516 29.776 28.26 ;
  LAYER M1 ;
        RECT 29.744 28.356 29.776 28.596 ;
  LAYER M1 ;
        RECT 29.744 28.692 29.776 29.436 ;
  LAYER M1 ;
        RECT 29.744 29.532 29.776 29.772 ;
  LAYER M1 ;
        RECT 29.744 29.868 29.776 30.612 ;
  LAYER M1 ;
        RECT 29.744 30.708 29.776 30.948 ;
  LAYER M1 ;
        RECT 29.744 31.044 29.776 31.788 ;
  LAYER M1 ;
        RECT 29.744 31.884 29.776 32.124 ;
  LAYER M1 ;
        RECT 29.744 32.22 29.776 32.964 ;
  LAYER M1 ;
        RECT 29.744 33.06 29.776 33.3 ;
  LAYER M1 ;
        RECT 29.744 33.396 29.776 34.14 ;
  LAYER M1 ;
        RECT 29.744 34.236 29.776 34.476 ;
  LAYER M1 ;
        RECT 29.744 34.572 29.776 35.316 ;
  LAYER M1 ;
        RECT 29.744 35.412 29.776 35.652 ;
  LAYER M1 ;
        RECT 29.744 35.748 29.776 36.492 ;
  LAYER M1 ;
        RECT 29.744 36.588 29.776 36.828 ;
  LAYER M1 ;
        RECT 29.744 37.092 29.776 37.332 ;
  LAYER M1 ;
        RECT 29.824 25.164 29.856 25.908 ;
  LAYER M1 ;
        RECT 29.824 26.34 29.856 27.084 ;
  LAYER M1 ;
        RECT 29.824 27.516 29.856 28.26 ;
  LAYER M1 ;
        RECT 29.824 28.692 29.856 29.436 ;
  LAYER M1 ;
        RECT 29.824 29.868 29.856 30.612 ;
  LAYER M1 ;
        RECT 29.824 31.044 29.856 31.788 ;
  LAYER M1 ;
        RECT 29.824 32.22 29.856 32.964 ;
  LAYER M1 ;
        RECT 29.824 33.396 29.856 34.14 ;
  LAYER M1 ;
        RECT 29.824 34.572 29.856 35.316 ;
  LAYER M1 ;
        RECT 29.824 35.748 29.856 36.492 ;
  LAYER M1 ;
        RECT 29.904 25.164 29.936 25.908 ;
  LAYER M1 ;
        RECT 29.904 26.004 29.936 26.244 ;
  LAYER M1 ;
        RECT 29.904 26.34 29.936 27.084 ;
  LAYER M1 ;
        RECT 29.904 27.18 29.936 27.42 ;
  LAYER M1 ;
        RECT 29.904 27.516 29.936 28.26 ;
  LAYER M1 ;
        RECT 29.904 28.356 29.936 28.596 ;
  LAYER M1 ;
        RECT 29.904 28.692 29.936 29.436 ;
  LAYER M1 ;
        RECT 29.904 29.532 29.936 29.772 ;
  LAYER M1 ;
        RECT 29.904 29.868 29.936 30.612 ;
  LAYER M1 ;
        RECT 29.904 30.708 29.936 30.948 ;
  LAYER M1 ;
        RECT 29.904 31.044 29.936 31.788 ;
  LAYER M1 ;
        RECT 29.904 31.884 29.936 32.124 ;
  LAYER M1 ;
        RECT 29.904 32.22 29.936 32.964 ;
  LAYER M1 ;
        RECT 29.904 33.06 29.936 33.3 ;
  LAYER M1 ;
        RECT 29.904 33.396 29.936 34.14 ;
  LAYER M1 ;
        RECT 29.904 34.236 29.936 34.476 ;
  LAYER M1 ;
        RECT 29.904 34.572 29.936 35.316 ;
  LAYER M1 ;
        RECT 29.904 35.412 29.936 35.652 ;
  LAYER M1 ;
        RECT 29.904 35.748 29.936 36.492 ;
  LAYER M1 ;
        RECT 29.904 36.588 29.936 36.828 ;
  LAYER M1 ;
        RECT 29.904 37.092 29.936 37.332 ;
  LAYER M1 ;
        RECT 29.984 25.164 30.016 25.908 ;
  LAYER M1 ;
        RECT 29.984 26.34 30.016 27.084 ;
  LAYER M1 ;
        RECT 29.984 27.516 30.016 28.26 ;
  LAYER M1 ;
        RECT 29.984 28.692 30.016 29.436 ;
  LAYER M1 ;
        RECT 29.984 29.868 30.016 30.612 ;
  LAYER M1 ;
        RECT 29.984 31.044 30.016 31.788 ;
  LAYER M1 ;
        RECT 29.984 32.22 30.016 32.964 ;
  LAYER M1 ;
        RECT 29.984 33.396 30.016 34.14 ;
  LAYER M1 ;
        RECT 29.984 34.572 30.016 35.316 ;
  LAYER M1 ;
        RECT 29.984 35.748 30.016 36.492 ;
  LAYER M1 ;
        RECT 30.064 25.164 30.096 25.908 ;
  LAYER M1 ;
        RECT 30.064 26.004 30.096 26.244 ;
  LAYER M1 ;
        RECT 30.064 26.34 30.096 27.084 ;
  LAYER M1 ;
        RECT 30.064 27.18 30.096 27.42 ;
  LAYER M1 ;
        RECT 30.064 27.516 30.096 28.26 ;
  LAYER M1 ;
        RECT 30.064 28.356 30.096 28.596 ;
  LAYER M1 ;
        RECT 30.064 28.692 30.096 29.436 ;
  LAYER M1 ;
        RECT 30.064 29.532 30.096 29.772 ;
  LAYER M1 ;
        RECT 30.064 29.868 30.096 30.612 ;
  LAYER M1 ;
        RECT 30.064 30.708 30.096 30.948 ;
  LAYER M1 ;
        RECT 30.064 31.044 30.096 31.788 ;
  LAYER M1 ;
        RECT 30.064 31.884 30.096 32.124 ;
  LAYER M1 ;
        RECT 30.064 32.22 30.096 32.964 ;
  LAYER M1 ;
        RECT 30.064 33.06 30.096 33.3 ;
  LAYER M1 ;
        RECT 30.064 33.396 30.096 34.14 ;
  LAYER M1 ;
        RECT 30.064 34.236 30.096 34.476 ;
  LAYER M1 ;
        RECT 30.064 34.572 30.096 35.316 ;
  LAYER M1 ;
        RECT 30.064 35.412 30.096 35.652 ;
  LAYER M1 ;
        RECT 30.064 35.748 30.096 36.492 ;
  LAYER M1 ;
        RECT 30.064 36.588 30.096 36.828 ;
  LAYER M1 ;
        RECT 30.064 37.092 30.096 37.332 ;
  LAYER M1 ;
        RECT 30.144 25.164 30.176 25.908 ;
  LAYER M1 ;
        RECT 30.144 26.34 30.176 27.084 ;
  LAYER M1 ;
        RECT 30.144 27.516 30.176 28.26 ;
  LAYER M1 ;
        RECT 30.144 28.692 30.176 29.436 ;
  LAYER M1 ;
        RECT 30.144 29.868 30.176 30.612 ;
  LAYER M1 ;
        RECT 30.144 31.044 30.176 31.788 ;
  LAYER M1 ;
        RECT 30.144 32.22 30.176 32.964 ;
  LAYER M1 ;
        RECT 30.144 33.396 30.176 34.14 ;
  LAYER M1 ;
        RECT 30.144 34.572 30.176 35.316 ;
  LAYER M1 ;
        RECT 30.144 35.748 30.176 36.492 ;
  LAYER M1 ;
        RECT 30.224 25.164 30.256 25.908 ;
  LAYER M1 ;
        RECT 30.224 26.004 30.256 26.244 ;
  LAYER M1 ;
        RECT 30.224 26.34 30.256 27.084 ;
  LAYER M1 ;
        RECT 30.224 27.18 30.256 27.42 ;
  LAYER M1 ;
        RECT 30.224 27.516 30.256 28.26 ;
  LAYER M1 ;
        RECT 30.224 28.356 30.256 28.596 ;
  LAYER M1 ;
        RECT 30.224 28.692 30.256 29.436 ;
  LAYER M1 ;
        RECT 30.224 29.532 30.256 29.772 ;
  LAYER M1 ;
        RECT 30.224 29.868 30.256 30.612 ;
  LAYER M1 ;
        RECT 30.224 30.708 30.256 30.948 ;
  LAYER M1 ;
        RECT 30.224 31.044 30.256 31.788 ;
  LAYER M1 ;
        RECT 30.224 31.884 30.256 32.124 ;
  LAYER M1 ;
        RECT 30.224 32.22 30.256 32.964 ;
  LAYER M1 ;
        RECT 30.224 33.06 30.256 33.3 ;
  LAYER M1 ;
        RECT 30.224 33.396 30.256 34.14 ;
  LAYER M1 ;
        RECT 30.224 34.236 30.256 34.476 ;
  LAYER M1 ;
        RECT 30.224 34.572 30.256 35.316 ;
  LAYER M1 ;
        RECT 30.224 35.412 30.256 35.652 ;
  LAYER M1 ;
        RECT 30.224 35.748 30.256 36.492 ;
  LAYER M1 ;
        RECT 30.224 36.588 30.256 36.828 ;
  LAYER M1 ;
        RECT 30.224 37.092 30.256 37.332 ;
  LAYER M1 ;
        RECT 30.304 25.164 30.336 25.908 ;
  LAYER M1 ;
        RECT 30.304 26.34 30.336 27.084 ;
  LAYER M1 ;
        RECT 30.304 27.516 30.336 28.26 ;
  LAYER M1 ;
        RECT 30.304 28.692 30.336 29.436 ;
  LAYER M1 ;
        RECT 30.304 29.868 30.336 30.612 ;
  LAYER M1 ;
        RECT 30.304 31.044 30.336 31.788 ;
  LAYER M1 ;
        RECT 30.304 32.22 30.336 32.964 ;
  LAYER M1 ;
        RECT 30.304 33.396 30.336 34.14 ;
  LAYER M1 ;
        RECT 30.304 34.572 30.336 35.316 ;
  LAYER M1 ;
        RECT 30.304 35.748 30.336 36.492 ;
  LAYER M1 ;
        RECT 30.384 25.164 30.416 25.908 ;
  LAYER M1 ;
        RECT 30.384 26.004 30.416 26.244 ;
  LAYER M1 ;
        RECT 30.384 26.34 30.416 27.084 ;
  LAYER M1 ;
        RECT 30.384 27.18 30.416 27.42 ;
  LAYER M1 ;
        RECT 30.384 27.516 30.416 28.26 ;
  LAYER M1 ;
        RECT 30.384 28.356 30.416 28.596 ;
  LAYER M1 ;
        RECT 30.384 28.692 30.416 29.436 ;
  LAYER M1 ;
        RECT 30.384 29.532 30.416 29.772 ;
  LAYER M1 ;
        RECT 30.384 29.868 30.416 30.612 ;
  LAYER M1 ;
        RECT 30.384 30.708 30.416 30.948 ;
  LAYER M1 ;
        RECT 30.384 31.044 30.416 31.788 ;
  LAYER M1 ;
        RECT 30.384 31.884 30.416 32.124 ;
  LAYER M1 ;
        RECT 30.384 32.22 30.416 32.964 ;
  LAYER M1 ;
        RECT 30.384 33.06 30.416 33.3 ;
  LAYER M1 ;
        RECT 30.384 33.396 30.416 34.14 ;
  LAYER M1 ;
        RECT 30.384 34.236 30.416 34.476 ;
  LAYER M1 ;
        RECT 30.384 34.572 30.416 35.316 ;
  LAYER M1 ;
        RECT 30.384 35.412 30.416 35.652 ;
  LAYER M1 ;
        RECT 30.384 35.748 30.416 36.492 ;
  LAYER M1 ;
        RECT 30.384 36.588 30.416 36.828 ;
  LAYER M1 ;
        RECT 30.384 37.092 30.416 37.332 ;
  LAYER M1 ;
        RECT 30.464 25.164 30.496 25.908 ;
  LAYER M1 ;
        RECT 30.464 26.34 30.496 27.084 ;
  LAYER M1 ;
        RECT 30.464 27.516 30.496 28.26 ;
  LAYER M1 ;
        RECT 30.464 28.692 30.496 29.436 ;
  LAYER M1 ;
        RECT 30.464 29.868 30.496 30.612 ;
  LAYER M1 ;
        RECT 30.464 31.044 30.496 31.788 ;
  LAYER M1 ;
        RECT 30.464 32.22 30.496 32.964 ;
  LAYER M1 ;
        RECT 30.464 33.396 30.496 34.14 ;
  LAYER M1 ;
        RECT 30.464 34.572 30.496 35.316 ;
  LAYER M1 ;
        RECT 30.464 35.748 30.496 36.492 ;
  LAYER M1 ;
        RECT 30.544 25.164 30.576 25.908 ;
  LAYER M1 ;
        RECT 30.544 26.004 30.576 26.244 ;
  LAYER M1 ;
        RECT 30.544 26.34 30.576 27.084 ;
  LAYER M1 ;
        RECT 30.544 27.18 30.576 27.42 ;
  LAYER M1 ;
        RECT 30.544 27.516 30.576 28.26 ;
  LAYER M1 ;
        RECT 30.544 28.356 30.576 28.596 ;
  LAYER M1 ;
        RECT 30.544 28.692 30.576 29.436 ;
  LAYER M1 ;
        RECT 30.544 29.532 30.576 29.772 ;
  LAYER M1 ;
        RECT 30.544 29.868 30.576 30.612 ;
  LAYER M1 ;
        RECT 30.544 30.708 30.576 30.948 ;
  LAYER M1 ;
        RECT 30.544 31.044 30.576 31.788 ;
  LAYER M1 ;
        RECT 30.544 31.884 30.576 32.124 ;
  LAYER M1 ;
        RECT 30.544 32.22 30.576 32.964 ;
  LAYER M1 ;
        RECT 30.544 33.06 30.576 33.3 ;
  LAYER M1 ;
        RECT 30.544 33.396 30.576 34.14 ;
  LAYER M1 ;
        RECT 30.544 34.236 30.576 34.476 ;
  LAYER M1 ;
        RECT 30.544 34.572 30.576 35.316 ;
  LAYER M1 ;
        RECT 30.544 35.412 30.576 35.652 ;
  LAYER M1 ;
        RECT 30.544 35.748 30.576 36.492 ;
  LAYER M1 ;
        RECT 30.544 36.588 30.576 36.828 ;
  LAYER M1 ;
        RECT 30.544 37.092 30.576 37.332 ;
  LAYER M1 ;
        RECT 30.624 25.164 30.656 25.908 ;
  LAYER M1 ;
        RECT 30.624 26.34 30.656 27.084 ;
  LAYER M1 ;
        RECT 30.624 27.516 30.656 28.26 ;
  LAYER M1 ;
        RECT 30.624 28.692 30.656 29.436 ;
  LAYER M1 ;
        RECT 30.624 29.868 30.656 30.612 ;
  LAYER M1 ;
        RECT 30.624 31.044 30.656 31.788 ;
  LAYER M1 ;
        RECT 30.624 32.22 30.656 32.964 ;
  LAYER M1 ;
        RECT 30.624 33.396 30.656 34.14 ;
  LAYER M1 ;
        RECT 30.624 34.572 30.656 35.316 ;
  LAYER M1 ;
        RECT 30.624 35.748 30.656 36.492 ;
  LAYER M1 ;
        RECT 30.704 25.164 30.736 25.908 ;
  LAYER M1 ;
        RECT 30.704 26.004 30.736 26.244 ;
  LAYER M1 ;
        RECT 30.704 26.34 30.736 27.084 ;
  LAYER M1 ;
        RECT 30.704 27.18 30.736 27.42 ;
  LAYER M1 ;
        RECT 30.704 27.516 30.736 28.26 ;
  LAYER M1 ;
        RECT 30.704 28.356 30.736 28.596 ;
  LAYER M1 ;
        RECT 30.704 28.692 30.736 29.436 ;
  LAYER M1 ;
        RECT 30.704 29.532 30.736 29.772 ;
  LAYER M1 ;
        RECT 30.704 29.868 30.736 30.612 ;
  LAYER M1 ;
        RECT 30.704 30.708 30.736 30.948 ;
  LAYER M1 ;
        RECT 30.704 31.044 30.736 31.788 ;
  LAYER M1 ;
        RECT 30.704 31.884 30.736 32.124 ;
  LAYER M1 ;
        RECT 30.704 32.22 30.736 32.964 ;
  LAYER M1 ;
        RECT 30.704 33.06 30.736 33.3 ;
  LAYER M1 ;
        RECT 30.704 33.396 30.736 34.14 ;
  LAYER M1 ;
        RECT 30.704 34.236 30.736 34.476 ;
  LAYER M1 ;
        RECT 30.704 34.572 30.736 35.316 ;
  LAYER M1 ;
        RECT 30.704 35.412 30.736 35.652 ;
  LAYER M1 ;
        RECT 30.704 35.748 30.736 36.492 ;
  LAYER M1 ;
        RECT 30.704 36.588 30.736 36.828 ;
  LAYER M1 ;
        RECT 30.704 37.092 30.736 37.332 ;
  LAYER M1 ;
        RECT 30.784 25.164 30.816 25.908 ;
  LAYER M1 ;
        RECT 30.784 26.34 30.816 27.084 ;
  LAYER M1 ;
        RECT 30.784 27.516 30.816 28.26 ;
  LAYER M1 ;
        RECT 30.784 28.692 30.816 29.436 ;
  LAYER M1 ;
        RECT 30.784 29.868 30.816 30.612 ;
  LAYER M1 ;
        RECT 30.784 31.044 30.816 31.788 ;
  LAYER M1 ;
        RECT 30.784 32.22 30.816 32.964 ;
  LAYER M1 ;
        RECT 30.784 33.396 30.816 34.14 ;
  LAYER M1 ;
        RECT 30.784 34.572 30.816 35.316 ;
  LAYER M1 ;
        RECT 30.784 35.748 30.816 36.492 ;
  LAYER M1 ;
        RECT 30.864 25.164 30.896 25.908 ;
  LAYER M1 ;
        RECT 30.864 26.004 30.896 26.244 ;
  LAYER M1 ;
        RECT 30.864 26.34 30.896 27.084 ;
  LAYER M1 ;
        RECT 30.864 27.18 30.896 27.42 ;
  LAYER M1 ;
        RECT 30.864 27.516 30.896 28.26 ;
  LAYER M1 ;
        RECT 30.864 28.356 30.896 28.596 ;
  LAYER M1 ;
        RECT 30.864 28.692 30.896 29.436 ;
  LAYER M1 ;
        RECT 30.864 29.532 30.896 29.772 ;
  LAYER M1 ;
        RECT 30.864 29.868 30.896 30.612 ;
  LAYER M1 ;
        RECT 30.864 30.708 30.896 30.948 ;
  LAYER M1 ;
        RECT 30.864 31.044 30.896 31.788 ;
  LAYER M1 ;
        RECT 30.864 31.884 30.896 32.124 ;
  LAYER M1 ;
        RECT 30.864 32.22 30.896 32.964 ;
  LAYER M1 ;
        RECT 30.864 33.06 30.896 33.3 ;
  LAYER M1 ;
        RECT 30.864 33.396 30.896 34.14 ;
  LAYER M1 ;
        RECT 30.864 34.236 30.896 34.476 ;
  LAYER M1 ;
        RECT 30.864 34.572 30.896 35.316 ;
  LAYER M1 ;
        RECT 30.864 35.412 30.896 35.652 ;
  LAYER M1 ;
        RECT 30.864 35.748 30.896 36.492 ;
  LAYER M1 ;
        RECT 30.864 36.588 30.896 36.828 ;
  LAYER M1 ;
        RECT 30.864 37.092 30.896 37.332 ;
  LAYER M1 ;
        RECT 30.944 25.164 30.976 25.908 ;
  LAYER M1 ;
        RECT 30.944 26.34 30.976 27.084 ;
  LAYER M1 ;
        RECT 30.944 27.516 30.976 28.26 ;
  LAYER M1 ;
        RECT 30.944 28.692 30.976 29.436 ;
  LAYER M1 ;
        RECT 30.944 29.868 30.976 30.612 ;
  LAYER M1 ;
        RECT 30.944 31.044 30.976 31.788 ;
  LAYER M1 ;
        RECT 30.944 32.22 30.976 32.964 ;
  LAYER M1 ;
        RECT 30.944 33.396 30.976 34.14 ;
  LAYER M1 ;
        RECT 30.944 34.572 30.976 35.316 ;
  LAYER M1 ;
        RECT 30.944 35.748 30.976 36.492 ;
  LAYER M1 ;
        RECT 31.024 25.164 31.056 25.908 ;
  LAYER M1 ;
        RECT 31.024 26.004 31.056 26.244 ;
  LAYER M1 ;
        RECT 31.024 26.34 31.056 27.084 ;
  LAYER M1 ;
        RECT 31.024 27.18 31.056 27.42 ;
  LAYER M1 ;
        RECT 31.024 27.516 31.056 28.26 ;
  LAYER M1 ;
        RECT 31.024 28.356 31.056 28.596 ;
  LAYER M1 ;
        RECT 31.024 28.692 31.056 29.436 ;
  LAYER M1 ;
        RECT 31.024 29.532 31.056 29.772 ;
  LAYER M1 ;
        RECT 31.024 29.868 31.056 30.612 ;
  LAYER M1 ;
        RECT 31.024 30.708 31.056 30.948 ;
  LAYER M1 ;
        RECT 31.024 31.044 31.056 31.788 ;
  LAYER M1 ;
        RECT 31.024 31.884 31.056 32.124 ;
  LAYER M1 ;
        RECT 31.024 32.22 31.056 32.964 ;
  LAYER M1 ;
        RECT 31.024 33.06 31.056 33.3 ;
  LAYER M1 ;
        RECT 31.024 33.396 31.056 34.14 ;
  LAYER M1 ;
        RECT 31.024 34.236 31.056 34.476 ;
  LAYER M1 ;
        RECT 31.024 34.572 31.056 35.316 ;
  LAYER M1 ;
        RECT 31.024 35.412 31.056 35.652 ;
  LAYER M1 ;
        RECT 31.024 35.748 31.056 36.492 ;
  LAYER M1 ;
        RECT 31.024 36.588 31.056 36.828 ;
  LAYER M1 ;
        RECT 31.024 37.092 31.056 37.332 ;
  LAYER M1 ;
        RECT 31.104 25.164 31.136 25.908 ;
  LAYER M1 ;
        RECT 31.104 26.34 31.136 27.084 ;
  LAYER M1 ;
        RECT 31.104 27.516 31.136 28.26 ;
  LAYER M1 ;
        RECT 31.104 28.692 31.136 29.436 ;
  LAYER M1 ;
        RECT 31.104 29.868 31.136 30.612 ;
  LAYER M1 ;
        RECT 31.104 31.044 31.136 31.788 ;
  LAYER M1 ;
        RECT 31.104 32.22 31.136 32.964 ;
  LAYER M1 ;
        RECT 31.104 33.396 31.136 34.14 ;
  LAYER M1 ;
        RECT 31.104 34.572 31.136 35.316 ;
  LAYER M1 ;
        RECT 31.104 35.748 31.136 36.492 ;
  LAYER M1 ;
        RECT 31.184 25.164 31.216 25.908 ;
  LAYER M1 ;
        RECT 31.184 26.004 31.216 26.244 ;
  LAYER M1 ;
        RECT 31.184 26.34 31.216 27.084 ;
  LAYER M1 ;
        RECT 31.184 27.18 31.216 27.42 ;
  LAYER M1 ;
        RECT 31.184 27.516 31.216 28.26 ;
  LAYER M1 ;
        RECT 31.184 28.356 31.216 28.596 ;
  LAYER M1 ;
        RECT 31.184 28.692 31.216 29.436 ;
  LAYER M1 ;
        RECT 31.184 29.532 31.216 29.772 ;
  LAYER M1 ;
        RECT 31.184 29.868 31.216 30.612 ;
  LAYER M1 ;
        RECT 31.184 30.708 31.216 30.948 ;
  LAYER M1 ;
        RECT 31.184 31.044 31.216 31.788 ;
  LAYER M1 ;
        RECT 31.184 31.884 31.216 32.124 ;
  LAYER M1 ;
        RECT 31.184 32.22 31.216 32.964 ;
  LAYER M1 ;
        RECT 31.184 33.06 31.216 33.3 ;
  LAYER M1 ;
        RECT 31.184 33.396 31.216 34.14 ;
  LAYER M1 ;
        RECT 31.184 34.236 31.216 34.476 ;
  LAYER M1 ;
        RECT 31.184 34.572 31.216 35.316 ;
  LAYER M1 ;
        RECT 31.184 35.412 31.216 35.652 ;
  LAYER M1 ;
        RECT 31.184 35.748 31.216 36.492 ;
  LAYER M1 ;
        RECT 31.184 36.588 31.216 36.828 ;
  LAYER M1 ;
        RECT 31.184 37.092 31.216 37.332 ;
  LAYER M1 ;
        RECT 31.264 25.164 31.296 25.908 ;
  LAYER M1 ;
        RECT 31.264 26.34 31.296 27.084 ;
  LAYER M1 ;
        RECT 31.264 27.516 31.296 28.26 ;
  LAYER M1 ;
        RECT 31.264 28.692 31.296 29.436 ;
  LAYER M1 ;
        RECT 31.264 29.868 31.296 30.612 ;
  LAYER M1 ;
        RECT 31.264 31.044 31.296 31.788 ;
  LAYER M1 ;
        RECT 31.264 32.22 31.296 32.964 ;
  LAYER M1 ;
        RECT 31.264 33.396 31.296 34.14 ;
  LAYER M1 ;
        RECT 31.264 34.572 31.296 35.316 ;
  LAYER M1 ;
        RECT 31.264 35.748 31.296 36.492 ;
  LAYER M1 ;
        RECT 31.344 25.164 31.376 25.908 ;
  LAYER M1 ;
        RECT 31.344 26.004 31.376 26.244 ;
  LAYER M1 ;
        RECT 31.344 26.34 31.376 27.084 ;
  LAYER M1 ;
        RECT 31.344 27.18 31.376 27.42 ;
  LAYER M1 ;
        RECT 31.344 27.516 31.376 28.26 ;
  LAYER M1 ;
        RECT 31.344 28.356 31.376 28.596 ;
  LAYER M1 ;
        RECT 31.344 28.692 31.376 29.436 ;
  LAYER M1 ;
        RECT 31.344 29.532 31.376 29.772 ;
  LAYER M1 ;
        RECT 31.344 29.868 31.376 30.612 ;
  LAYER M1 ;
        RECT 31.344 30.708 31.376 30.948 ;
  LAYER M1 ;
        RECT 31.344 31.044 31.376 31.788 ;
  LAYER M1 ;
        RECT 31.344 31.884 31.376 32.124 ;
  LAYER M1 ;
        RECT 31.344 32.22 31.376 32.964 ;
  LAYER M1 ;
        RECT 31.344 33.06 31.376 33.3 ;
  LAYER M1 ;
        RECT 31.344 33.396 31.376 34.14 ;
  LAYER M1 ;
        RECT 31.344 34.236 31.376 34.476 ;
  LAYER M1 ;
        RECT 31.344 34.572 31.376 35.316 ;
  LAYER M1 ;
        RECT 31.344 35.412 31.376 35.652 ;
  LAYER M1 ;
        RECT 31.344 35.748 31.376 36.492 ;
  LAYER M1 ;
        RECT 31.344 36.588 31.376 36.828 ;
  LAYER M1 ;
        RECT 31.344 37.092 31.376 37.332 ;
  LAYER M1 ;
        RECT 31.424 25.164 31.456 25.908 ;
  LAYER M1 ;
        RECT 31.424 26.34 31.456 27.084 ;
  LAYER M1 ;
        RECT 31.424 27.516 31.456 28.26 ;
  LAYER M1 ;
        RECT 31.424 28.692 31.456 29.436 ;
  LAYER M1 ;
        RECT 31.424 29.868 31.456 30.612 ;
  LAYER M1 ;
        RECT 31.424 31.044 31.456 31.788 ;
  LAYER M1 ;
        RECT 31.424 32.22 31.456 32.964 ;
  LAYER M1 ;
        RECT 31.424 33.396 31.456 34.14 ;
  LAYER M1 ;
        RECT 31.424 34.572 31.456 35.316 ;
  LAYER M1 ;
        RECT 31.424 35.748 31.456 36.492 ;
  LAYER M1 ;
        RECT 31.504 25.164 31.536 25.908 ;
  LAYER M1 ;
        RECT 31.504 26.004 31.536 26.244 ;
  LAYER M1 ;
        RECT 31.504 26.34 31.536 27.084 ;
  LAYER M1 ;
        RECT 31.504 27.18 31.536 27.42 ;
  LAYER M1 ;
        RECT 31.504 27.516 31.536 28.26 ;
  LAYER M1 ;
        RECT 31.504 28.356 31.536 28.596 ;
  LAYER M1 ;
        RECT 31.504 28.692 31.536 29.436 ;
  LAYER M1 ;
        RECT 31.504 29.532 31.536 29.772 ;
  LAYER M1 ;
        RECT 31.504 29.868 31.536 30.612 ;
  LAYER M1 ;
        RECT 31.504 30.708 31.536 30.948 ;
  LAYER M1 ;
        RECT 31.504 31.044 31.536 31.788 ;
  LAYER M1 ;
        RECT 31.504 31.884 31.536 32.124 ;
  LAYER M1 ;
        RECT 31.504 32.22 31.536 32.964 ;
  LAYER M1 ;
        RECT 31.504 33.06 31.536 33.3 ;
  LAYER M1 ;
        RECT 31.504 33.396 31.536 34.14 ;
  LAYER M1 ;
        RECT 31.504 34.236 31.536 34.476 ;
  LAYER M1 ;
        RECT 31.504 34.572 31.536 35.316 ;
  LAYER M1 ;
        RECT 31.504 35.412 31.536 35.652 ;
  LAYER M1 ;
        RECT 31.504 35.748 31.536 36.492 ;
  LAYER M1 ;
        RECT 31.504 36.588 31.536 36.828 ;
  LAYER M1 ;
        RECT 31.504 37.092 31.536 37.332 ;
  LAYER M1 ;
        RECT 31.584 25.164 31.616 25.908 ;
  LAYER M1 ;
        RECT 31.584 26.34 31.616 27.084 ;
  LAYER M1 ;
        RECT 31.584 27.516 31.616 28.26 ;
  LAYER M1 ;
        RECT 31.584 28.692 31.616 29.436 ;
  LAYER M1 ;
        RECT 31.584 29.868 31.616 30.612 ;
  LAYER M1 ;
        RECT 31.584 31.044 31.616 31.788 ;
  LAYER M1 ;
        RECT 31.584 32.22 31.616 32.964 ;
  LAYER M1 ;
        RECT 31.584 33.396 31.616 34.14 ;
  LAYER M1 ;
        RECT 31.584 34.572 31.616 35.316 ;
  LAYER M1 ;
        RECT 31.584 35.748 31.616 36.492 ;
  LAYER M2 ;
        RECT 27.564 25.184 31.636 25.216 ;
  LAYER M2 ;
        RECT 27.644 25.268 31.556 25.3 ;
  LAYER M2 ;
        RECT 27.644 26.024 31.556 26.056 ;
  LAYER M2 ;
        RECT 27.564 26.36 31.636 26.392 ;
  LAYER M2 ;
        RECT 27.644 26.444 31.556 26.476 ;
  LAYER M2 ;
        RECT 27.644 27.2 31.556 27.232 ;
  LAYER M2 ;
        RECT 27.564 27.536 31.636 27.568 ;
  LAYER M2 ;
        RECT 27.644 27.62 31.556 27.652 ;
  LAYER M2 ;
        RECT 27.644 28.376 31.556 28.408 ;
  LAYER M2 ;
        RECT 27.564 28.712 31.636 28.744 ;
  LAYER M2 ;
        RECT 27.644 28.796 31.556 28.828 ;
  LAYER M2 ;
        RECT 27.644 29.552 31.556 29.584 ;
  LAYER M2 ;
        RECT 27.564 29.888 31.636 29.92 ;
  LAYER M2 ;
        RECT 27.644 29.972 31.556 30.004 ;
  LAYER M2 ;
        RECT 27.644 30.728 31.556 30.76 ;
  LAYER M2 ;
        RECT 27.564 31.064 31.636 31.096 ;
  LAYER M2 ;
        RECT 27.644 31.148 31.556 31.18 ;
  LAYER M2 ;
        RECT 27.644 31.904 31.556 31.936 ;
  LAYER M2 ;
        RECT 27.564 32.24 31.636 32.272 ;
  LAYER M2 ;
        RECT 27.644 32.324 31.556 32.356 ;
  LAYER M2 ;
        RECT 27.644 33.08 31.556 33.112 ;
  LAYER M2 ;
        RECT 27.564 33.416 31.636 33.448 ;
  LAYER M2 ;
        RECT 27.644 33.5 31.556 33.532 ;
  LAYER M2 ;
        RECT 27.644 34.256 31.556 34.288 ;
  LAYER M2 ;
        RECT 27.564 34.592 31.636 34.624 ;
  LAYER M2 ;
        RECT 27.644 34.676 31.556 34.708 ;
  LAYER M2 ;
        RECT 27.644 35.432 31.556 35.464 ;
  LAYER M2 ;
        RECT 27.564 35.768 31.636 35.8 ;
  LAYER M2 ;
        RECT 27.644 35.852 31.556 35.884 ;
  LAYER M2 ;
        RECT 27.644 36.608 31.556 36.64 ;
  LAYER M1 ;
        RECT 5.184 9.372 5.216 15.576 ;
  LAYER M1 ;
        RECT 5.184 15.524 5.28 15.556 ;
  LAYER M1 ;
        RECT 5.248 9.372 5.28 15.576 ;
  LAYER M1 ;
        RECT 5.248 9.392 5.344 9.424 ;
  LAYER M1 ;
        RECT 5.312 9.372 5.344 15.576 ;
  LAYER M1 ;
        RECT 5.312 15.524 5.408 15.556 ;
  LAYER M1 ;
        RECT 5.376 9.372 5.408 15.576 ;
  LAYER M1 ;
        RECT 5.376 9.392 5.472 9.424 ;
  LAYER M1 ;
        RECT 5.44 9.372 5.472 15.576 ;
  LAYER M1 ;
        RECT 5.44 15.524 5.536 15.556 ;
  LAYER M1 ;
        RECT 5.504 9.372 5.536 15.576 ;
  LAYER M1 ;
        RECT 5.504 9.392 5.6 9.424 ;
  LAYER M1 ;
        RECT 5.568 9.372 5.6 15.576 ;
  LAYER M1 ;
        RECT 5.568 15.524 5.664 15.556 ;
  LAYER M1 ;
        RECT 5.632 9.372 5.664 15.576 ;
  LAYER M1 ;
        RECT 5.632 9.392 5.728 9.424 ;
  LAYER M1 ;
        RECT 5.696 9.372 5.728 15.576 ;
  LAYER M1 ;
        RECT 5.696 15.524 5.792 15.556 ;
  LAYER M1 ;
        RECT 5.76 9.372 5.792 15.576 ;
  LAYER M1 ;
        RECT 5.76 9.392 5.856 9.424 ;
  LAYER M1 ;
        RECT 5.824 9.372 5.856 15.576 ;
  LAYER M1 ;
        RECT 5.824 15.524 5.92 15.556 ;
  LAYER M1 ;
        RECT 5.888 9.372 5.92 15.576 ;
  LAYER M1 ;
        RECT 5.888 9.392 5.984 9.424 ;
  LAYER M1 ;
        RECT 5.952 9.372 5.984 15.576 ;
  LAYER M1 ;
        RECT 5.952 15.524 6.048 15.556 ;
  LAYER M1 ;
        RECT 6.016 9.372 6.048 15.576 ;
  LAYER M1 ;
        RECT 6.016 9.392 6.112 9.424 ;
  LAYER M1 ;
        RECT 6.08 9.372 6.112 15.576 ;
  LAYER M1 ;
        RECT 6.08 15.524 6.176 15.556 ;
  LAYER M1 ;
        RECT 6.144 9.372 6.176 15.576 ;
  LAYER M1 ;
        RECT 6.144 9.392 6.24 9.424 ;
  LAYER M1 ;
        RECT 6.208 9.372 6.24 15.576 ;
  LAYER M1 ;
        RECT 6.208 15.524 6.304 15.556 ;
  LAYER M1 ;
        RECT 6.272 9.372 6.304 15.576 ;
  LAYER M1 ;
        RECT 6.272 9.392 6.368 9.424 ;
  LAYER M1 ;
        RECT 6.336 9.372 6.368 15.576 ;
  LAYER M1 ;
        RECT 6.336 15.524 6.432 15.556 ;
  LAYER M1 ;
        RECT 6.4 9.372 6.432 15.576 ;
  LAYER M1 ;
        RECT 6.4 9.392 6.496 9.424 ;
  LAYER M1 ;
        RECT 6.464 9.372 6.496 15.576 ;
  LAYER M1 ;
        RECT 6.464 15.524 6.56 15.556 ;
  LAYER M1 ;
        RECT 6.528 9.372 6.56 15.576 ;
  LAYER M1 ;
        RECT 0.064 0.048 0.096 18.348 ;
  LAYER M1 ;
        RECT 0.064 18.296 0.16 18.328 ;
  LAYER M1 ;
        RECT 0.128 0.048 0.16 18.348 ;
  LAYER M1 ;
        RECT 0.128 0.068 0.224 0.1 ;
  LAYER M1 ;
        RECT 0.192 0.048 0.224 18.348 ;
  LAYER M1 ;
        RECT 0.192 18.296 0.288 18.328 ;
  LAYER M1 ;
        RECT 0.256 0.048 0.288 18.348 ;
  LAYER M1 ;
        RECT 0.256 0.068 0.352 0.1 ;
  LAYER M1 ;
        RECT 0.32 0.048 0.352 18.348 ;
  LAYER M1 ;
        RECT 0.32 18.296 0.416 18.328 ;
  LAYER M1 ;
        RECT 0.384 0.048 0.416 18.348 ;
  LAYER M1 ;
        RECT 0.384 0.068 0.48 0.1 ;
  LAYER M1 ;
        RECT 0.448 0.048 0.48 18.348 ;
  LAYER M1 ;
        RECT 0.448 18.296 0.544 18.328 ;
  LAYER M1 ;
        RECT 0.512 0.048 0.544 18.348 ;
  LAYER M1 ;
        RECT 0.512 0.068 0.608 0.1 ;
  LAYER M1 ;
        RECT 0.576 0.048 0.608 18.348 ;
  LAYER M1 ;
        RECT 0.576 18.296 0.672 18.328 ;
  LAYER M1 ;
        RECT 0.64 0.048 0.672 18.348 ;
  LAYER M1 ;
        RECT 0.64 0.068 0.736 0.1 ;
  LAYER M1 ;
        RECT 0.704 0.048 0.736 18.348 ;
  LAYER M1 ;
        RECT 0.704 18.296 0.8 18.328 ;
  LAYER M1 ;
        RECT 0.768 0.048 0.8 18.348 ;
  LAYER M1 ;
        RECT 0.768 0.068 0.864 0.1 ;
  LAYER M1 ;
        RECT 0.832 0.048 0.864 18.348 ;
  LAYER M1 ;
        RECT 0.832 18.296 0.928 18.328 ;
  LAYER M1 ;
        RECT 0.896 0.048 0.928 18.348 ;
  LAYER M1 ;
        RECT 0.896 0.068 0.992 0.1 ;
  LAYER M1 ;
        RECT 0.96 0.048 0.992 18.348 ;
  LAYER M1 ;
        RECT 0.96 18.296 1.056 18.328 ;
  LAYER M1 ;
        RECT 1.024 0.048 1.056 18.348 ;
  LAYER M1 ;
        RECT 1.024 0.068 1.12 0.1 ;
  LAYER M1 ;
        RECT 1.088 0.048 1.12 18.348 ;
  LAYER M1 ;
        RECT 1.088 18.296 1.184 18.328 ;
  LAYER M1 ;
        RECT 1.152 0.048 1.184 18.348 ;
  LAYER M1 ;
        RECT 1.152 0.068 1.248 0.1 ;
  LAYER M1 ;
        RECT 1.216 0.048 1.248 18.348 ;
  LAYER M1 ;
        RECT 1.216 18.296 1.312 18.328 ;
  LAYER M1 ;
        RECT 1.28 0.048 1.312 18.348 ;
  LAYER M1 ;
        RECT 1.28 0.068 1.376 0.1 ;
  LAYER M1 ;
        RECT 1.344 0.048 1.376 18.348 ;
  LAYER M1 ;
        RECT 1.344 18.296 1.44 18.328 ;
  LAYER M1 ;
        RECT 1.408 0.048 1.44 18.348 ;
  LAYER M1 ;
        RECT 1.408 0.068 1.504 0.1 ;
  LAYER M1 ;
        RECT 1.472 0.048 1.504 18.348 ;
  LAYER M1 ;
        RECT 1.472 18.296 1.568 18.328 ;
  LAYER M1 ;
        RECT 1.536 0.048 1.568 18.348 ;
  LAYER M1 ;
        RECT 1.536 0.068 1.632 0.1 ;
  LAYER M1 ;
        RECT 1.6 0.048 1.632 18.348 ;
  LAYER M1 ;
        RECT 1.6 18.296 1.696 18.328 ;
  LAYER M1 ;
        RECT 1.664 0.048 1.696 18.348 ;
  LAYER M1 ;
        RECT 1.664 0.068 1.76 0.1 ;
  LAYER M1 ;
        RECT 1.728 0.048 1.76 18.348 ;
  LAYER M1 ;
        RECT 1.728 18.296 1.824 18.328 ;
  LAYER M1 ;
        RECT 1.792 0.048 1.824 18.348 ;
  LAYER M1 ;
        RECT 1.792 0.068 1.888 0.1 ;
  LAYER M1 ;
        RECT 1.856 0.048 1.888 18.348 ;
  LAYER M1 ;
        RECT 1.856 18.296 1.952 18.328 ;
  LAYER M1 ;
        RECT 1.92 0.048 1.952 18.348 ;
  LAYER M1 ;
        RECT 1.92 0.068 2.016 0.1 ;
  LAYER M1 ;
        RECT 1.984 0.048 2.016 18.348 ;
  LAYER M1 ;
        RECT 1.984 18.296 2.08 18.328 ;
  LAYER M1 ;
        RECT 2.048 0.048 2.08 18.348 ;
  LAYER M1 ;
        RECT 2.048 0.068 2.144 0.1 ;
  LAYER M1 ;
        RECT 2.112 0.048 2.144 18.348 ;
  LAYER M1 ;
        RECT 2.112 18.296 2.208 18.328 ;
  LAYER M1 ;
        RECT 2.176 0.048 2.208 18.348 ;
  LAYER M1 ;
        RECT 2.176 0.068 2.272 0.1 ;
  LAYER M1 ;
        RECT 2.24 0.048 2.272 18.348 ;
  LAYER M1 ;
        RECT 2.24 18.296 2.336 18.328 ;
  LAYER M1 ;
        RECT 2.304 0.048 2.336 18.348 ;
  LAYER M1 ;
        RECT 2.304 0.068 2.4 0.1 ;
  LAYER M1 ;
        RECT 2.368 0.048 2.4 18.348 ;
  LAYER M1 ;
        RECT 2.368 18.296 2.464 18.328 ;
  LAYER M1 ;
        RECT 2.432 0.048 2.464 18.348 ;
  LAYER M1 ;
        RECT 2.432 0.068 2.528 0.1 ;
  LAYER M1 ;
        RECT 2.496 0.048 2.528 18.348 ;
  LAYER M1 ;
        RECT 2.496 18.296 2.592 18.328 ;
  LAYER M1 ;
        RECT 2.56 0.048 2.592 18.348 ;
  LAYER M1 ;
        RECT 2.56 0.068 2.656 0.1 ;
  LAYER M1 ;
        RECT 2.624 0.048 2.656 18.348 ;
  LAYER M1 ;
        RECT 2.624 18.296 2.72 18.328 ;
  LAYER M1 ;
        RECT 2.688 0.048 2.72 18.348 ;
  LAYER M1 ;
        RECT 2.688 0.068 2.784 0.1 ;
  LAYER M1 ;
        RECT 2.752 0.048 2.784 18.348 ;
  LAYER M1 ;
        RECT 2.752 18.296 2.848 18.328 ;
  LAYER M1 ;
        RECT 2.816 0.048 2.848 18.348 ;
  LAYER M1 ;
        RECT 2.816 0.068 2.912 0.1 ;
  LAYER M1 ;
        RECT 2.88 0.048 2.912 18.348 ;
  LAYER M1 ;
        RECT 2.88 18.296 2.976 18.328 ;
  LAYER M1 ;
        RECT 2.944 0.048 2.976 18.348 ;
  LAYER M1 ;
        RECT 2.944 0.068 3.04 0.1 ;
  LAYER M1 ;
        RECT 3.008 0.048 3.04 18.348 ;
  LAYER M1 ;
        RECT 3.008 18.296 3.104 18.328 ;
  LAYER M1 ;
        RECT 3.072 0.048 3.104 18.348 ;
  LAYER M1 ;
        RECT 3.072 0.068 3.168 0.1 ;
  LAYER M1 ;
        RECT 3.136 0.048 3.168 18.348 ;
  LAYER M1 ;
        RECT 3.136 18.296 3.232 18.328 ;
  LAYER M1 ;
        RECT 3.2 0.048 3.232 18.348 ;
  LAYER M1 ;
        RECT 3.2 0.068 3.296 0.1 ;
  LAYER M1 ;
        RECT 3.264 0.048 3.296 18.348 ;
  LAYER M1 ;
        RECT 3.264 18.296 3.36 18.328 ;
  LAYER M1 ;
        RECT 3.328 0.048 3.36 18.348 ;
  LAYER M1 ;
        RECT 3.328 0.068 3.424 0.1 ;
  LAYER M1 ;
        RECT 3.392 0.048 3.424 18.348 ;
  LAYER M1 ;
        RECT 3.392 18.296 3.488 18.328 ;
  LAYER M1 ;
        RECT 3.456 0.048 3.488 18.348 ;
  LAYER M1 ;
        RECT 3.456 0.068 3.552 0.1 ;
  LAYER M1 ;
        RECT 3.52 0.048 3.552 18.348 ;
  LAYER M1 ;
        RECT 3.52 18.296 3.616 18.328 ;
  LAYER M1 ;
        RECT 3.584 0.048 3.616 18.348 ;
  LAYER M1 ;
        RECT 3.584 0.068 3.68 0.1 ;
  LAYER M1 ;
        RECT 3.648 0.048 3.68 18.348 ;
  LAYER M1 ;
        RECT 3.648 18.296 3.744 18.328 ;
  LAYER M1 ;
        RECT 3.712 0.048 3.744 18.348 ;
  LAYER M1 ;
        RECT 3.712 0.068 3.808 0.1 ;
  LAYER M1 ;
        RECT 3.776 0.048 3.808 18.348 ;
  LAYER M1 ;
        RECT 3.776 18.296 3.872 18.328 ;
  LAYER M1 ;
        RECT 3.84 0.048 3.872 18.348 ;
  LAYER M1 ;
        RECT 3.84 0.068 3.936 0.1 ;
  LAYER M1 ;
        RECT 3.904 0.048 3.936 18.348 ;
  LAYER M1 ;
        RECT 3.904 18.296 4 18.328 ;
  LAYER M1 ;
        RECT 3.968 0.048 4 18.348 ;
  LAYER M1 ;
        RECT 3.968 0.068 4.064 0.1 ;
  LAYER M1 ;
        RECT 4.032 0.048 4.064 18.348 ;
  LAYER M1 ;
        RECT 11.664 0.216 11.696 0.96 ;
  LAYER M1 ;
        RECT 11.664 1.056 11.696 1.296 ;
  LAYER M1 ;
        RECT 11.664 1.392 11.696 2.136 ;
  LAYER M1 ;
        RECT 11.664 2.232 11.696 2.472 ;
  LAYER M1 ;
        RECT 11.664 2.568 11.696 3.312 ;
  LAYER M1 ;
        RECT 11.664 3.408 11.696 3.648 ;
  LAYER M1 ;
        RECT 11.664 3.744 11.696 4.488 ;
  LAYER M1 ;
        RECT 11.664 4.584 11.696 4.824 ;
  LAYER M1 ;
        RECT 11.664 4.92 11.696 5.664 ;
  LAYER M1 ;
        RECT 11.664 5.76 11.696 6 ;
  LAYER M1 ;
        RECT 11.664 6.096 11.696 6.84 ;
  LAYER M1 ;
        RECT 11.664 6.936 11.696 7.176 ;
  LAYER M1 ;
        RECT 11.664 7.272 11.696 8.016 ;
  LAYER M1 ;
        RECT 11.664 8.112 11.696 8.352 ;
  LAYER M1 ;
        RECT 11.664 8.616 11.696 8.856 ;
  LAYER M1 ;
        RECT 11.584 0.216 11.616 0.96 ;
  LAYER M1 ;
        RECT 11.584 1.392 11.616 2.136 ;
  LAYER M1 ;
        RECT 11.584 2.568 11.616 3.312 ;
  LAYER M1 ;
        RECT 11.584 3.744 11.616 4.488 ;
  LAYER M1 ;
        RECT 11.584 4.92 11.616 5.664 ;
  LAYER M1 ;
        RECT 11.584 6.096 11.616 6.84 ;
  LAYER M1 ;
        RECT 11.584 7.272 11.616 8.016 ;
  LAYER M1 ;
        RECT 11.744 0.216 11.776 0.96 ;
  LAYER M1 ;
        RECT 11.744 1.392 11.776 2.136 ;
  LAYER M1 ;
        RECT 11.744 2.568 11.776 3.312 ;
  LAYER M1 ;
        RECT 11.744 3.744 11.776 4.488 ;
  LAYER M1 ;
        RECT 11.744 4.92 11.776 5.664 ;
  LAYER M1 ;
        RECT 11.744 6.096 11.776 6.84 ;
  LAYER M1 ;
        RECT 11.744 7.272 11.776 8.016 ;
  LAYER M1 ;
        RECT 11.824 0.216 11.856 0.96 ;
  LAYER M1 ;
        RECT 11.824 1.056 11.856 1.296 ;
  LAYER M1 ;
        RECT 11.824 1.392 11.856 2.136 ;
  LAYER M1 ;
        RECT 11.824 2.232 11.856 2.472 ;
  LAYER M1 ;
        RECT 11.824 2.568 11.856 3.312 ;
  LAYER M1 ;
        RECT 11.824 3.408 11.856 3.648 ;
  LAYER M1 ;
        RECT 11.824 3.744 11.856 4.488 ;
  LAYER M1 ;
        RECT 11.824 4.584 11.856 4.824 ;
  LAYER M1 ;
        RECT 11.824 4.92 11.856 5.664 ;
  LAYER M1 ;
        RECT 11.824 5.76 11.856 6 ;
  LAYER M1 ;
        RECT 11.824 6.096 11.856 6.84 ;
  LAYER M1 ;
        RECT 11.824 6.936 11.856 7.176 ;
  LAYER M1 ;
        RECT 11.824 7.272 11.856 8.016 ;
  LAYER M1 ;
        RECT 11.824 8.112 11.856 8.352 ;
  LAYER M1 ;
        RECT 11.824 8.616 11.856 8.856 ;
  LAYER M1 ;
        RECT 11.904 0.216 11.936 0.96 ;
  LAYER M1 ;
        RECT 11.904 1.392 11.936 2.136 ;
  LAYER M1 ;
        RECT 11.904 2.568 11.936 3.312 ;
  LAYER M1 ;
        RECT 11.904 3.744 11.936 4.488 ;
  LAYER M1 ;
        RECT 11.904 4.92 11.936 5.664 ;
  LAYER M1 ;
        RECT 11.904 6.096 11.936 6.84 ;
  LAYER M1 ;
        RECT 11.904 7.272 11.936 8.016 ;
  LAYER M1 ;
        RECT 11.984 0.216 12.016 0.96 ;
  LAYER M1 ;
        RECT 11.984 1.056 12.016 1.296 ;
  LAYER M1 ;
        RECT 11.984 1.392 12.016 2.136 ;
  LAYER M1 ;
        RECT 11.984 2.232 12.016 2.472 ;
  LAYER M1 ;
        RECT 11.984 2.568 12.016 3.312 ;
  LAYER M1 ;
        RECT 11.984 3.408 12.016 3.648 ;
  LAYER M1 ;
        RECT 11.984 3.744 12.016 4.488 ;
  LAYER M1 ;
        RECT 11.984 4.584 12.016 4.824 ;
  LAYER M1 ;
        RECT 11.984 4.92 12.016 5.664 ;
  LAYER M1 ;
        RECT 11.984 5.76 12.016 6 ;
  LAYER M1 ;
        RECT 11.984 6.096 12.016 6.84 ;
  LAYER M1 ;
        RECT 11.984 6.936 12.016 7.176 ;
  LAYER M1 ;
        RECT 11.984 7.272 12.016 8.016 ;
  LAYER M1 ;
        RECT 11.984 8.112 12.016 8.352 ;
  LAYER M1 ;
        RECT 11.984 8.616 12.016 8.856 ;
  LAYER M1 ;
        RECT 12.064 0.216 12.096 0.96 ;
  LAYER M1 ;
        RECT 12.064 1.392 12.096 2.136 ;
  LAYER M1 ;
        RECT 12.064 2.568 12.096 3.312 ;
  LAYER M1 ;
        RECT 12.064 3.744 12.096 4.488 ;
  LAYER M1 ;
        RECT 12.064 4.92 12.096 5.664 ;
  LAYER M1 ;
        RECT 12.064 6.096 12.096 6.84 ;
  LAYER M1 ;
        RECT 12.064 7.272 12.096 8.016 ;
  LAYER M1 ;
        RECT 12.144 0.216 12.176 0.96 ;
  LAYER M1 ;
        RECT 12.144 1.056 12.176 1.296 ;
  LAYER M1 ;
        RECT 12.144 1.392 12.176 2.136 ;
  LAYER M1 ;
        RECT 12.144 2.232 12.176 2.472 ;
  LAYER M1 ;
        RECT 12.144 2.568 12.176 3.312 ;
  LAYER M1 ;
        RECT 12.144 3.408 12.176 3.648 ;
  LAYER M1 ;
        RECT 12.144 3.744 12.176 4.488 ;
  LAYER M1 ;
        RECT 12.144 4.584 12.176 4.824 ;
  LAYER M1 ;
        RECT 12.144 4.92 12.176 5.664 ;
  LAYER M1 ;
        RECT 12.144 5.76 12.176 6 ;
  LAYER M1 ;
        RECT 12.144 6.096 12.176 6.84 ;
  LAYER M1 ;
        RECT 12.144 6.936 12.176 7.176 ;
  LAYER M1 ;
        RECT 12.144 7.272 12.176 8.016 ;
  LAYER M1 ;
        RECT 12.144 8.112 12.176 8.352 ;
  LAYER M1 ;
        RECT 12.144 8.616 12.176 8.856 ;
  LAYER M1 ;
        RECT 12.224 0.216 12.256 0.96 ;
  LAYER M1 ;
        RECT 12.224 1.392 12.256 2.136 ;
  LAYER M1 ;
        RECT 12.224 2.568 12.256 3.312 ;
  LAYER M1 ;
        RECT 12.224 3.744 12.256 4.488 ;
  LAYER M1 ;
        RECT 12.224 4.92 12.256 5.664 ;
  LAYER M1 ;
        RECT 12.224 6.096 12.256 6.84 ;
  LAYER M1 ;
        RECT 12.224 7.272 12.256 8.016 ;
  LAYER M1 ;
        RECT 12.304 0.216 12.336 0.96 ;
  LAYER M1 ;
        RECT 12.304 1.056 12.336 1.296 ;
  LAYER M1 ;
        RECT 12.304 1.392 12.336 2.136 ;
  LAYER M1 ;
        RECT 12.304 2.232 12.336 2.472 ;
  LAYER M1 ;
        RECT 12.304 2.568 12.336 3.312 ;
  LAYER M1 ;
        RECT 12.304 3.408 12.336 3.648 ;
  LAYER M1 ;
        RECT 12.304 3.744 12.336 4.488 ;
  LAYER M1 ;
        RECT 12.304 4.584 12.336 4.824 ;
  LAYER M1 ;
        RECT 12.304 4.92 12.336 5.664 ;
  LAYER M1 ;
        RECT 12.304 5.76 12.336 6 ;
  LAYER M1 ;
        RECT 12.304 6.096 12.336 6.84 ;
  LAYER M1 ;
        RECT 12.304 6.936 12.336 7.176 ;
  LAYER M1 ;
        RECT 12.304 7.272 12.336 8.016 ;
  LAYER M1 ;
        RECT 12.304 8.112 12.336 8.352 ;
  LAYER M1 ;
        RECT 12.304 8.616 12.336 8.856 ;
  LAYER M1 ;
        RECT 12.384 0.216 12.416 0.96 ;
  LAYER M1 ;
        RECT 12.384 1.392 12.416 2.136 ;
  LAYER M1 ;
        RECT 12.384 2.568 12.416 3.312 ;
  LAYER M1 ;
        RECT 12.384 3.744 12.416 4.488 ;
  LAYER M1 ;
        RECT 12.384 4.92 12.416 5.664 ;
  LAYER M1 ;
        RECT 12.384 6.096 12.416 6.84 ;
  LAYER M1 ;
        RECT 12.384 7.272 12.416 8.016 ;
  LAYER M1 ;
        RECT 12.464 0.216 12.496 0.96 ;
  LAYER M1 ;
        RECT 12.464 1.056 12.496 1.296 ;
  LAYER M1 ;
        RECT 12.464 1.392 12.496 2.136 ;
  LAYER M1 ;
        RECT 12.464 2.232 12.496 2.472 ;
  LAYER M1 ;
        RECT 12.464 2.568 12.496 3.312 ;
  LAYER M1 ;
        RECT 12.464 3.408 12.496 3.648 ;
  LAYER M1 ;
        RECT 12.464 3.744 12.496 4.488 ;
  LAYER M1 ;
        RECT 12.464 4.584 12.496 4.824 ;
  LAYER M1 ;
        RECT 12.464 4.92 12.496 5.664 ;
  LAYER M1 ;
        RECT 12.464 5.76 12.496 6 ;
  LAYER M1 ;
        RECT 12.464 6.096 12.496 6.84 ;
  LAYER M1 ;
        RECT 12.464 6.936 12.496 7.176 ;
  LAYER M1 ;
        RECT 12.464 7.272 12.496 8.016 ;
  LAYER M1 ;
        RECT 12.464 8.112 12.496 8.352 ;
  LAYER M1 ;
        RECT 12.464 8.616 12.496 8.856 ;
  LAYER M1 ;
        RECT 12.544 0.216 12.576 0.96 ;
  LAYER M1 ;
        RECT 12.544 1.392 12.576 2.136 ;
  LAYER M1 ;
        RECT 12.544 2.568 12.576 3.312 ;
  LAYER M1 ;
        RECT 12.544 3.744 12.576 4.488 ;
  LAYER M1 ;
        RECT 12.544 4.92 12.576 5.664 ;
  LAYER M1 ;
        RECT 12.544 6.096 12.576 6.84 ;
  LAYER M1 ;
        RECT 12.544 7.272 12.576 8.016 ;
  LAYER M1 ;
        RECT 12.624 0.216 12.656 0.96 ;
  LAYER M1 ;
        RECT 12.624 1.056 12.656 1.296 ;
  LAYER M1 ;
        RECT 12.624 1.392 12.656 2.136 ;
  LAYER M1 ;
        RECT 12.624 2.232 12.656 2.472 ;
  LAYER M1 ;
        RECT 12.624 2.568 12.656 3.312 ;
  LAYER M1 ;
        RECT 12.624 3.408 12.656 3.648 ;
  LAYER M1 ;
        RECT 12.624 3.744 12.656 4.488 ;
  LAYER M1 ;
        RECT 12.624 4.584 12.656 4.824 ;
  LAYER M1 ;
        RECT 12.624 4.92 12.656 5.664 ;
  LAYER M1 ;
        RECT 12.624 5.76 12.656 6 ;
  LAYER M1 ;
        RECT 12.624 6.096 12.656 6.84 ;
  LAYER M1 ;
        RECT 12.624 6.936 12.656 7.176 ;
  LAYER M1 ;
        RECT 12.624 7.272 12.656 8.016 ;
  LAYER M1 ;
        RECT 12.624 8.112 12.656 8.352 ;
  LAYER M1 ;
        RECT 12.624 8.616 12.656 8.856 ;
  LAYER M1 ;
        RECT 12.704 0.216 12.736 0.96 ;
  LAYER M1 ;
        RECT 12.704 1.392 12.736 2.136 ;
  LAYER M1 ;
        RECT 12.704 2.568 12.736 3.312 ;
  LAYER M1 ;
        RECT 12.704 3.744 12.736 4.488 ;
  LAYER M1 ;
        RECT 12.704 4.92 12.736 5.664 ;
  LAYER M1 ;
        RECT 12.704 6.096 12.736 6.84 ;
  LAYER M1 ;
        RECT 12.704 7.272 12.736 8.016 ;
  LAYER M1 ;
        RECT 12.784 0.216 12.816 0.96 ;
  LAYER M1 ;
        RECT 12.784 1.056 12.816 1.296 ;
  LAYER M1 ;
        RECT 12.784 1.392 12.816 2.136 ;
  LAYER M1 ;
        RECT 12.784 2.232 12.816 2.472 ;
  LAYER M1 ;
        RECT 12.784 2.568 12.816 3.312 ;
  LAYER M1 ;
        RECT 12.784 3.408 12.816 3.648 ;
  LAYER M1 ;
        RECT 12.784 3.744 12.816 4.488 ;
  LAYER M1 ;
        RECT 12.784 4.584 12.816 4.824 ;
  LAYER M1 ;
        RECT 12.784 4.92 12.816 5.664 ;
  LAYER M1 ;
        RECT 12.784 5.76 12.816 6 ;
  LAYER M1 ;
        RECT 12.784 6.096 12.816 6.84 ;
  LAYER M1 ;
        RECT 12.784 6.936 12.816 7.176 ;
  LAYER M1 ;
        RECT 12.784 7.272 12.816 8.016 ;
  LAYER M1 ;
        RECT 12.784 8.112 12.816 8.352 ;
  LAYER M1 ;
        RECT 12.784 8.616 12.816 8.856 ;
  LAYER M1 ;
        RECT 12.864 0.216 12.896 0.96 ;
  LAYER M1 ;
        RECT 12.864 1.392 12.896 2.136 ;
  LAYER M1 ;
        RECT 12.864 2.568 12.896 3.312 ;
  LAYER M1 ;
        RECT 12.864 3.744 12.896 4.488 ;
  LAYER M1 ;
        RECT 12.864 4.92 12.896 5.664 ;
  LAYER M1 ;
        RECT 12.864 6.096 12.896 6.84 ;
  LAYER M1 ;
        RECT 12.864 7.272 12.896 8.016 ;
  LAYER M1 ;
        RECT 12.944 0.216 12.976 0.96 ;
  LAYER M1 ;
        RECT 12.944 1.056 12.976 1.296 ;
  LAYER M1 ;
        RECT 12.944 1.392 12.976 2.136 ;
  LAYER M1 ;
        RECT 12.944 2.232 12.976 2.472 ;
  LAYER M1 ;
        RECT 12.944 2.568 12.976 3.312 ;
  LAYER M1 ;
        RECT 12.944 3.408 12.976 3.648 ;
  LAYER M1 ;
        RECT 12.944 3.744 12.976 4.488 ;
  LAYER M1 ;
        RECT 12.944 4.584 12.976 4.824 ;
  LAYER M1 ;
        RECT 12.944 4.92 12.976 5.664 ;
  LAYER M1 ;
        RECT 12.944 5.76 12.976 6 ;
  LAYER M1 ;
        RECT 12.944 6.096 12.976 6.84 ;
  LAYER M1 ;
        RECT 12.944 6.936 12.976 7.176 ;
  LAYER M1 ;
        RECT 12.944 7.272 12.976 8.016 ;
  LAYER M1 ;
        RECT 12.944 8.112 12.976 8.352 ;
  LAYER M1 ;
        RECT 12.944 8.616 12.976 8.856 ;
  LAYER M1 ;
        RECT 13.024 0.216 13.056 0.96 ;
  LAYER M1 ;
        RECT 13.024 1.392 13.056 2.136 ;
  LAYER M1 ;
        RECT 13.024 2.568 13.056 3.312 ;
  LAYER M1 ;
        RECT 13.024 3.744 13.056 4.488 ;
  LAYER M1 ;
        RECT 13.024 4.92 13.056 5.664 ;
  LAYER M1 ;
        RECT 13.024 6.096 13.056 6.84 ;
  LAYER M1 ;
        RECT 13.024 7.272 13.056 8.016 ;
  LAYER M1 ;
        RECT 13.104 0.216 13.136 0.96 ;
  LAYER M1 ;
        RECT 13.104 1.056 13.136 1.296 ;
  LAYER M1 ;
        RECT 13.104 1.392 13.136 2.136 ;
  LAYER M1 ;
        RECT 13.104 2.232 13.136 2.472 ;
  LAYER M1 ;
        RECT 13.104 2.568 13.136 3.312 ;
  LAYER M1 ;
        RECT 13.104 3.408 13.136 3.648 ;
  LAYER M1 ;
        RECT 13.104 3.744 13.136 4.488 ;
  LAYER M1 ;
        RECT 13.104 4.584 13.136 4.824 ;
  LAYER M1 ;
        RECT 13.104 4.92 13.136 5.664 ;
  LAYER M1 ;
        RECT 13.104 5.76 13.136 6 ;
  LAYER M1 ;
        RECT 13.104 6.096 13.136 6.84 ;
  LAYER M1 ;
        RECT 13.104 6.936 13.136 7.176 ;
  LAYER M1 ;
        RECT 13.104 7.272 13.136 8.016 ;
  LAYER M1 ;
        RECT 13.104 8.112 13.136 8.352 ;
  LAYER M1 ;
        RECT 13.104 8.616 13.136 8.856 ;
  LAYER M1 ;
        RECT 13.184 0.216 13.216 0.96 ;
  LAYER M1 ;
        RECT 13.184 1.392 13.216 2.136 ;
  LAYER M1 ;
        RECT 13.184 2.568 13.216 3.312 ;
  LAYER M1 ;
        RECT 13.184 3.744 13.216 4.488 ;
  LAYER M1 ;
        RECT 13.184 4.92 13.216 5.664 ;
  LAYER M1 ;
        RECT 13.184 6.096 13.216 6.84 ;
  LAYER M1 ;
        RECT 13.184 7.272 13.216 8.016 ;
  LAYER M1 ;
        RECT 13.264 0.216 13.296 0.96 ;
  LAYER M1 ;
        RECT 13.264 1.056 13.296 1.296 ;
  LAYER M1 ;
        RECT 13.264 1.392 13.296 2.136 ;
  LAYER M1 ;
        RECT 13.264 2.232 13.296 2.472 ;
  LAYER M1 ;
        RECT 13.264 2.568 13.296 3.312 ;
  LAYER M1 ;
        RECT 13.264 3.408 13.296 3.648 ;
  LAYER M1 ;
        RECT 13.264 3.744 13.296 4.488 ;
  LAYER M1 ;
        RECT 13.264 4.584 13.296 4.824 ;
  LAYER M1 ;
        RECT 13.264 4.92 13.296 5.664 ;
  LAYER M1 ;
        RECT 13.264 5.76 13.296 6 ;
  LAYER M1 ;
        RECT 13.264 6.096 13.296 6.84 ;
  LAYER M1 ;
        RECT 13.264 6.936 13.296 7.176 ;
  LAYER M1 ;
        RECT 13.264 7.272 13.296 8.016 ;
  LAYER M1 ;
        RECT 13.264 8.112 13.296 8.352 ;
  LAYER M1 ;
        RECT 13.264 8.616 13.296 8.856 ;
  LAYER M1 ;
        RECT 13.344 0.216 13.376 0.96 ;
  LAYER M1 ;
        RECT 13.344 1.392 13.376 2.136 ;
  LAYER M1 ;
        RECT 13.344 2.568 13.376 3.312 ;
  LAYER M1 ;
        RECT 13.344 3.744 13.376 4.488 ;
  LAYER M1 ;
        RECT 13.344 4.92 13.376 5.664 ;
  LAYER M1 ;
        RECT 13.344 6.096 13.376 6.84 ;
  LAYER M1 ;
        RECT 13.344 7.272 13.376 8.016 ;
  LAYER M1 ;
        RECT 13.424 0.216 13.456 0.96 ;
  LAYER M1 ;
        RECT 13.424 1.056 13.456 1.296 ;
  LAYER M1 ;
        RECT 13.424 1.392 13.456 2.136 ;
  LAYER M1 ;
        RECT 13.424 2.232 13.456 2.472 ;
  LAYER M1 ;
        RECT 13.424 2.568 13.456 3.312 ;
  LAYER M1 ;
        RECT 13.424 3.408 13.456 3.648 ;
  LAYER M1 ;
        RECT 13.424 3.744 13.456 4.488 ;
  LAYER M1 ;
        RECT 13.424 4.584 13.456 4.824 ;
  LAYER M1 ;
        RECT 13.424 4.92 13.456 5.664 ;
  LAYER M1 ;
        RECT 13.424 5.76 13.456 6 ;
  LAYER M1 ;
        RECT 13.424 6.096 13.456 6.84 ;
  LAYER M1 ;
        RECT 13.424 6.936 13.456 7.176 ;
  LAYER M1 ;
        RECT 13.424 7.272 13.456 8.016 ;
  LAYER M1 ;
        RECT 13.424 8.112 13.456 8.352 ;
  LAYER M1 ;
        RECT 13.424 8.616 13.456 8.856 ;
  LAYER M1 ;
        RECT 13.504 0.216 13.536 0.96 ;
  LAYER M1 ;
        RECT 13.504 1.392 13.536 2.136 ;
  LAYER M1 ;
        RECT 13.504 2.568 13.536 3.312 ;
  LAYER M1 ;
        RECT 13.504 3.744 13.536 4.488 ;
  LAYER M1 ;
        RECT 13.504 4.92 13.536 5.664 ;
  LAYER M1 ;
        RECT 13.504 6.096 13.536 6.84 ;
  LAYER M1 ;
        RECT 13.504 7.272 13.536 8.016 ;
  LAYER M2 ;
        RECT 11.564 0.236 13.556 0.268 ;
  LAYER M2 ;
        RECT 11.644 0.32 13.476 0.352 ;
  LAYER M2 ;
        RECT 11.644 1.076 13.476 1.108 ;
  LAYER M2 ;
        RECT 11.564 1.412 13.556 1.444 ;
  LAYER M2 ;
        RECT 11.644 1.496 13.476 1.528 ;
  LAYER M2 ;
        RECT 11.644 2.252 13.476 2.284 ;
  LAYER M2 ;
        RECT 11.564 2.588 13.556 2.62 ;
  LAYER M2 ;
        RECT 11.644 2.672 13.476 2.704 ;
  LAYER M2 ;
        RECT 11.644 3.428 13.476 3.46 ;
  LAYER M2 ;
        RECT 11.564 3.764 13.556 3.796 ;
  LAYER M2 ;
        RECT 11.644 3.848 13.476 3.88 ;
  LAYER M2 ;
        RECT 11.644 4.604 13.476 4.636 ;
  LAYER M2 ;
        RECT 11.564 4.94 13.556 4.972 ;
  LAYER M2 ;
        RECT 11.644 5.024 13.476 5.056 ;
  LAYER M2 ;
        RECT 11.644 5.78 13.476 5.812 ;
  LAYER M2 ;
        RECT 11.564 6.116 13.556 6.148 ;
  LAYER M2 ;
        RECT 11.644 6.2 13.476 6.232 ;
  LAYER M2 ;
        RECT 11.644 6.956 13.476 6.988 ;
  LAYER M2 ;
        RECT 11.564 7.292 13.556 7.324 ;
  LAYER M2 ;
        RECT 11.644 7.376 13.476 7.408 ;
  LAYER M2 ;
        RECT 11.644 8.132 13.476 8.164 ;
  LAYER M1 ;
        RECT 14.224 0.3 14.256 1.044 ;
  LAYER M1 ;
        RECT 14.224 1.14 14.256 1.38 ;
  LAYER M1 ;
        RECT 14.224 1.476 14.256 2.22 ;
  LAYER M1 ;
        RECT 14.224 2.316 14.256 2.556 ;
  LAYER M1 ;
        RECT 14.224 2.652 14.256 3.396 ;
  LAYER M1 ;
        RECT 14.224 3.492 14.256 3.732 ;
  LAYER M1 ;
        RECT 14.224 3.828 14.256 4.572 ;
  LAYER M1 ;
        RECT 14.224 4.668 14.256 4.908 ;
  LAYER M1 ;
        RECT 14.224 5.004 14.256 5.748 ;
  LAYER M1 ;
        RECT 14.224 5.844 14.256 6.084 ;
  LAYER M1 ;
        RECT 14.224 6.18 14.256 6.924 ;
  LAYER M1 ;
        RECT 14.224 7.02 14.256 7.26 ;
  LAYER M1 ;
        RECT 14.224 7.356 14.256 8.1 ;
  LAYER M1 ;
        RECT 14.224 8.196 14.256 8.436 ;
  LAYER M1 ;
        RECT 14.224 8.7 14.256 8.94 ;
  LAYER M1 ;
        RECT 14.144 0.3 14.176 1.044 ;
  LAYER M1 ;
        RECT 14.144 1.476 14.176 2.22 ;
  LAYER M1 ;
        RECT 14.144 2.652 14.176 3.396 ;
  LAYER M1 ;
        RECT 14.144 3.828 14.176 4.572 ;
  LAYER M1 ;
        RECT 14.144 5.004 14.176 5.748 ;
  LAYER M1 ;
        RECT 14.144 6.18 14.176 6.924 ;
  LAYER M1 ;
        RECT 14.144 7.356 14.176 8.1 ;
  LAYER M1 ;
        RECT 14.304 0.3 14.336 1.044 ;
  LAYER M1 ;
        RECT 14.304 1.476 14.336 2.22 ;
  LAYER M1 ;
        RECT 14.304 2.652 14.336 3.396 ;
  LAYER M1 ;
        RECT 14.304 3.828 14.336 4.572 ;
  LAYER M1 ;
        RECT 14.304 5.004 14.336 5.748 ;
  LAYER M1 ;
        RECT 14.304 6.18 14.336 6.924 ;
  LAYER M1 ;
        RECT 14.304 7.356 14.336 8.1 ;
  LAYER M1 ;
        RECT 14.384 0.3 14.416 1.044 ;
  LAYER M1 ;
        RECT 14.384 1.14 14.416 1.38 ;
  LAYER M1 ;
        RECT 14.384 1.476 14.416 2.22 ;
  LAYER M1 ;
        RECT 14.384 2.316 14.416 2.556 ;
  LAYER M1 ;
        RECT 14.384 2.652 14.416 3.396 ;
  LAYER M1 ;
        RECT 14.384 3.492 14.416 3.732 ;
  LAYER M1 ;
        RECT 14.384 3.828 14.416 4.572 ;
  LAYER M1 ;
        RECT 14.384 4.668 14.416 4.908 ;
  LAYER M1 ;
        RECT 14.384 5.004 14.416 5.748 ;
  LAYER M1 ;
        RECT 14.384 5.844 14.416 6.084 ;
  LAYER M1 ;
        RECT 14.384 6.18 14.416 6.924 ;
  LAYER M1 ;
        RECT 14.384 7.02 14.416 7.26 ;
  LAYER M1 ;
        RECT 14.384 7.356 14.416 8.1 ;
  LAYER M1 ;
        RECT 14.384 8.196 14.416 8.436 ;
  LAYER M1 ;
        RECT 14.384 8.7 14.416 8.94 ;
  LAYER M1 ;
        RECT 14.464 0.3 14.496 1.044 ;
  LAYER M1 ;
        RECT 14.464 1.476 14.496 2.22 ;
  LAYER M1 ;
        RECT 14.464 2.652 14.496 3.396 ;
  LAYER M1 ;
        RECT 14.464 3.828 14.496 4.572 ;
  LAYER M1 ;
        RECT 14.464 5.004 14.496 5.748 ;
  LAYER M1 ;
        RECT 14.464 6.18 14.496 6.924 ;
  LAYER M1 ;
        RECT 14.464 7.356 14.496 8.1 ;
  LAYER M1 ;
        RECT 14.544 0.3 14.576 1.044 ;
  LAYER M1 ;
        RECT 14.544 1.14 14.576 1.38 ;
  LAYER M1 ;
        RECT 14.544 1.476 14.576 2.22 ;
  LAYER M1 ;
        RECT 14.544 2.316 14.576 2.556 ;
  LAYER M1 ;
        RECT 14.544 2.652 14.576 3.396 ;
  LAYER M1 ;
        RECT 14.544 3.492 14.576 3.732 ;
  LAYER M1 ;
        RECT 14.544 3.828 14.576 4.572 ;
  LAYER M1 ;
        RECT 14.544 4.668 14.576 4.908 ;
  LAYER M1 ;
        RECT 14.544 5.004 14.576 5.748 ;
  LAYER M1 ;
        RECT 14.544 5.844 14.576 6.084 ;
  LAYER M1 ;
        RECT 14.544 6.18 14.576 6.924 ;
  LAYER M1 ;
        RECT 14.544 7.02 14.576 7.26 ;
  LAYER M1 ;
        RECT 14.544 7.356 14.576 8.1 ;
  LAYER M1 ;
        RECT 14.544 8.196 14.576 8.436 ;
  LAYER M1 ;
        RECT 14.544 8.7 14.576 8.94 ;
  LAYER M1 ;
        RECT 14.624 0.3 14.656 1.044 ;
  LAYER M1 ;
        RECT 14.624 1.476 14.656 2.22 ;
  LAYER M1 ;
        RECT 14.624 2.652 14.656 3.396 ;
  LAYER M1 ;
        RECT 14.624 3.828 14.656 4.572 ;
  LAYER M1 ;
        RECT 14.624 5.004 14.656 5.748 ;
  LAYER M1 ;
        RECT 14.624 6.18 14.656 6.924 ;
  LAYER M1 ;
        RECT 14.624 7.356 14.656 8.1 ;
  LAYER M1 ;
        RECT 14.704 0.3 14.736 1.044 ;
  LAYER M1 ;
        RECT 14.704 1.14 14.736 1.38 ;
  LAYER M1 ;
        RECT 14.704 1.476 14.736 2.22 ;
  LAYER M1 ;
        RECT 14.704 2.316 14.736 2.556 ;
  LAYER M1 ;
        RECT 14.704 2.652 14.736 3.396 ;
  LAYER M1 ;
        RECT 14.704 3.492 14.736 3.732 ;
  LAYER M1 ;
        RECT 14.704 3.828 14.736 4.572 ;
  LAYER M1 ;
        RECT 14.704 4.668 14.736 4.908 ;
  LAYER M1 ;
        RECT 14.704 5.004 14.736 5.748 ;
  LAYER M1 ;
        RECT 14.704 5.844 14.736 6.084 ;
  LAYER M1 ;
        RECT 14.704 6.18 14.736 6.924 ;
  LAYER M1 ;
        RECT 14.704 7.02 14.736 7.26 ;
  LAYER M1 ;
        RECT 14.704 7.356 14.736 8.1 ;
  LAYER M1 ;
        RECT 14.704 8.196 14.736 8.436 ;
  LAYER M1 ;
        RECT 14.704 8.7 14.736 8.94 ;
  LAYER M1 ;
        RECT 14.784 0.3 14.816 1.044 ;
  LAYER M1 ;
        RECT 14.784 1.476 14.816 2.22 ;
  LAYER M1 ;
        RECT 14.784 2.652 14.816 3.396 ;
  LAYER M1 ;
        RECT 14.784 3.828 14.816 4.572 ;
  LAYER M1 ;
        RECT 14.784 5.004 14.816 5.748 ;
  LAYER M1 ;
        RECT 14.784 6.18 14.816 6.924 ;
  LAYER M1 ;
        RECT 14.784 7.356 14.816 8.1 ;
  LAYER M1 ;
        RECT 14.864 0.3 14.896 1.044 ;
  LAYER M1 ;
        RECT 14.864 1.14 14.896 1.38 ;
  LAYER M1 ;
        RECT 14.864 1.476 14.896 2.22 ;
  LAYER M1 ;
        RECT 14.864 2.316 14.896 2.556 ;
  LAYER M1 ;
        RECT 14.864 2.652 14.896 3.396 ;
  LAYER M1 ;
        RECT 14.864 3.492 14.896 3.732 ;
  LAYER M1 ;
        RECT 14.864 3.828 14.896 4.572 ;
  LAYER M1 ;
        RECT 14.864 4.668 14.896 4.908 ;
  LAYER M1 ;
        RECT 14.864 5.004 14.896 5.748 ;
  LAYER M1 ;
        RECT 14.864 5.844 14.896 6.084 ;
  LAYER M1 ;
        RECT 14.864 6.18 14.896 6.924 ;
  LAYER M1 ;
        RECT 14.864 7.02 14.896 7.26 ;
  LAYER M1 ;
        RECT 14.864 7.356 14.896 8.1 ;
  LAYER M1 ;
        RECT 14.864 8.196 14.896 8.436 ;
  LAYER M1 ;
        RECT 14.864 8.7 14.896 8.94 ;
  LAYER M1 ;
        RECT 14.944 0.3 14.976 1.044 ;
  LAYER M1 ;
        RECT 14.944 1.476 14.976 2.22 ;
  LAYER M1 ;
        RECT 14.944 2.652 14.976 3.396 ;
  LAYER M1 ;
        RECT 14.944 3.828 14.976 4.572 ;
  LAYER M1 ;
        RECT 14.944 5.004 14.976 5.748 ;
  LAYER M1 ;
        RECT 14.944 6.18 14.976 6.924 ;
  LAYER M1 ;
        RECT 14.944 7.356 14.976 8.1 ;
  LAYER M1 ;
        RECT 15.024 0.3 15.056 1.044 ;
  LAYER M1 ;
        RECT 15.024 1.14 15.056 1.38 ;
  LAYER M1 ;
        RECT 15.024 1.476 15.056 2.22 ;
  LAYER M1 ;
        RECT 15.024 2.316 15.056 2.556 ;
  LAYER M1 ;
        RECT 15.024 2.652 15.056 3.396 ;
  LAYER M1 ;
        RECT 15.024 3.492 15.056 3.732 ;
  LAYER M1 ;
        RECT 15.024 3.828 15.056 4.572 ;
  LAYER M1 ;
        RECT 15.024 4.668 15.056 4.908 ;
  LAYER M1 ;
        RECT 15.024 5.004 15.056 5.748 ;
  LAYER M1 ;
        RECT 15.024 5.844 15.056 6.084 ;
  LAYER M1 ;
        RECT 15.024 6.18 15.056 6.924 ;
  LAYER M1 ;
        RECT 15.024 7.02 15.056 7.26 ;
  LAYER M1 ;
        RECT 15.024 7.356 15.056 8.1 ;
  LAYER M1 ;
        RECT 15.024 8.196 15.056 8.436 ;
  LAYER M1 ;
        RECT 15.024 8.7 15.056 8.94 ;
  LAYER M1 ;
        RECT 15.104 0.3 15.136 1.044 ;
  LAYER M1 ;
        RECT 15.104 1.476 15.136 2.22 ;
  LAYER M1 ;
        RECT 15.104 2.652 15.136 3.396 ;
  LAYER M1 ;
        RECT 15.104 3.828 15.136 4.572 ;
  LAYER M1 ;
        RECT 15.104 5.004 15.136 5.748 ;
  LAYER M1 ;
        RECT 15.104 6.18 15.136 6.924 ;
  LAYER M1 ;
        RECT 15.104 7.356 15.136 8.1 ;
  LAYER M1 ;
        RECT 15.184 0.3 15.216 1.044 ;
  LAYER M1 ;
        RECT 15.184 1.14 15.216 1.38 ;
  LAYER M1 ;
        RECT 15.184 1.476 15.216 2.22 ;
  LAYER M1 ;
        RECT 15.184 2.316 15.216 2.556 ;
  LAYER M1 ;
        RECT 15.184 2.652 15.216 3.396 ;
  LAYER M1 ;
        RECT 15.184 3.492 15.216 3.732 ;
  LAYER M1 ;
        RECT 15.184 3.828 15.216 4.572 ;
  LAYER M1 ;
        RECT 15.184 4.668 15.216 4.908 ;
  LAYER M1 ;
        RECT 15.184 5.004 15.216 5.748 ;
  LAYER M1 ;
        RECT 15.184 5.844 15.216 6.084 ;
  LAYER M1 ;
        RECT 15.184 6.18 15.216 6.924 ;
  LAYER M1 ;
        RECT 15.184 7.02 15.216 7.26 ;
  LAYER M1 ;
        RECT 15.184 7.356 15.216 8.1 ;
  LAYER M1 ;
        RECT 15.184 8.196 15.216 8.436 ;
  LAYER M1 ;
        RECT 15.184 8.7 15.216 8.94 ;
  LAYER M1 ;
        RECT 15.264 0.3 15.296 1.044 ;
  LAYER M1 ;
        RECT 15.264 1.476 15.296 2.22 ;
  LAYER M1 ;
        RECT 15.264 2.652 15.296 3.396 ;
  LAYER M1 ;
        RECT 15.264 3.828 15.296 4.572 ;
  LAYER M1 ;
        RECT 15.264 5.004 15.296 5.748 ;
  LAYER M1 ;
        RECT 15.264 6.18 15.296 6.924 ;
  LAYER M1 ;
        RECT 15.264 7.356 15.296 8.1 ;
  LAYER M1 ;
        RECT 15.344 0.3 15.376 1.044 ;
  LAYER M1 ;
        RECT 15.344 1.14 15.376 1.38 ;
  LAYER M1 ;
        RECT 15.344 1.476 15.376 2.22 ;
  LAYER M1 ;
        RECT 15.344 2.316 15.376 2.556 ;
  LAYER M1 ;
        RECT 15.344 2.652 15.376 3.396 ;
  LAYER M1 ;
        RECT 15.344 3.492 15.376 3.732 ;
  LAYER M1 ;
        RECT 15.344 3.828 15.376 4.572 ;
  LAYER M1 ;
        RECT 15.344 4.668 15.376 4.908 ;
  LAYER M1 ;
        RECT 15.344 5.004 15.376 5.748 ;
  LAYER M1 ;
        RECT 15.344 5.844 15.376 6.084 ;
  LAYER M1 ;
        RECT 15.344 6.18 15.376 6.924 ;
  LAYER M1 ;
        RECT 15.344 7.02 15.376 7.26 ;
  LAYER M1 ;
        RECT 15.344 7.356 15.376 8.1 ;
  LAYER M1 ;
        RECT 15.344 8.196 15.376 8.436 ;
  LAYER M1 ;
        RECT 15.344 8.7 15.376 8.94 ;
  LAYER M1 ;
        RECT 15.424 0.3 15.456 1.044 ;
  LAYER M1 ;
        RECT 15.424 1.476 15.456 2.22 ;
  LAYER M1 ;
        RECT 15.424 2.652 15.456 3.396 ;
  LAYER M1 ;
        RECT 15.424 3.828 15.456 4.572 ;
  LAYER M1 ;
        RECT 15.424 5.004 15.456 5.748 ;
  LAYER M1 ;
        RECT 15.424 6.18 15.456 6.924 ;
  LAYER M1 ;
        RECT 15.424 7.356 15.456 8.1 ;
  LAYER M1 ;
        RECT 15.504 0.3 15.536 1.044 ;
  LAYER M1 ;
        RECT 15.504 1.14 15.536 1.38 ;
  LAYER M1 ;
        RECT 15.504 1.476 15.536 2.22 ;
  LAYER M1 ;
        RECT 15.504 2.316 15.536 2.556 ;
  LAYER M1 ;
        RECT 15.504 2.652 15.536 3.396 ;
  LAYER M1 ;
        RECT 15.504 3.492 15.536 3.732 ;
  LAYER M1 ;
        RECT 15.504 3.828 15.536 4.572 ;
  LAYER M1 ;
        RECT 15.504 4.668 15.536 4.908 ;
  LAYER M1 ;
        RECT 15.504 5.004 15.536 5.748 ;
  LAYER M1 ;
        RECT 15.504 5.844 15.536 6.084 ;
  LAYER M1 ;
        RECT 15.504 6.18 15.536 6.924 ;
  LAYER M1 ;
        RECT 15.504 7.02 15.536 7.26 ;
  LAYER M1 ;
        RECT 15.504 7.356 15.536 8.1 ;
  LAYER M1 ;
        RECT 15.504 8.196 15.536 8.436 ;
  LAYER M1 ;
        RECT 15.504 8.7 15.536 8.94 ;
  LAYER M1 ;
        RECT 15.584 0.3 15.616 1.044 ;
  LAYER M1 ;
        RECT 15.584 1.476 15.616 2.22 ;
  LAYER M1 ;
        RECT 15.584 2.652 15.616 3.396 ;
  LAYER M1 ;
        RECT 15.584 3.828 15.616 4.572 ;
  LAYER M1 ;
        RECT 15.584 5.004 15.616 5.748 ;
  LAYER M1 ;
        RECT 15.584 6.18 15.616 6.924 ;
  LAYER M1 ;
        RECT 15.584 7.356 15.616 8.1 ;
  LAYER M1 ;
        RECT 15.664 0.3 15.696 1.044 ;
  LAYER M1 ;
        RECT 15.664 1.14 15.696 1.38 ;
  LAYER M1 ;
        RECT 15.664 1.476 15.696 2.22 ;
  LAYER M1 ;
        RECT 15.664 2.316 15.696 2.556 ;
  LAYER M1 ;
        RECT 15.664 2.652 15.696 3.396 ;
  LAYER M1 ;
        RECT 15.664 3.492 15.696 3.732 ;
  LAYER M1 ;
        RECT 15.664 3.828 15.696 4.572 ;
  LAYER M1 ;
        RECT 15.664 4.668 15.696 4.908 ;
  LAYER M1 ;
        RECT 15.664 5.004 15.696 5.748 ;
  LAYER M1 ;
        RECT 15.664 5.844 15.696 6.084 ;
  LAYER M1 ;
        RECT 15.664 6.18 15.696 6.924 ;
  LAYER M1 ;
        RECT 15.664 7.02 15.696 7.26 ;
  LAYER M1 ;
        RECT 15.664 7.356 15.696 8.1 ;
  LAYER M1 ;
        RECT 15.664 8.196 15.696 8.436 ;
  LAYER M1 ;
        RECT 15.664 8.7 15.696 8.94 ;
  LAYER M1 ;
        RECT 15.744 0.3 15.776 1.044 ;
  LAYER M1 ;
        RECT 15.744 1.476 15.776 2.22 ;
  LAYER M1 ;
        RECT 15.744 2.652 15.776 3.396 ;
  LAYER M1 ;
        RECT 15.744 3.828 15.776 4.572 ;
  LAYER M1 ;
        RECT 15.744 5.004 15.776 5.748 ;
  LAYER M1 ;
        RECT 15.744 6.18 15.776 6.924 ;
  LAYER M1 ;
        RECT 15.744 7.356 15.776 8.1 ;
  LAYER M1 ;
        RECT 15.824 0.3 15.856 1.044 ;
  LAYER M1 ;
        RECT 15.824 1.14 15.856 1.38 ;
  LAYER M1 ;
        RECT 15.824 1.476 15.856 2.22 ;
  LAYER M1 ;
        RECT 15.824 2.316 15.856 2.556 ;
  LAYER M1 ;
        RECT 15.824 2.652 15.856 3.396 ;
  LAYER M1 ;
        RECT 15.824 3.492 15.856 3.732 ;
  LAYER M1 ;
        RECT 15.824 3.828 15.856 4.572 ;
  LAYER M1 ;
        RECT 15.824 4.668 15.856 4.908 ;
  LAYER M1 ;
        RECT 15.824 5.004 15.856 5.748 ;
  LAYER M1 ;
        RECT 15.824 5.844 15.856 6.084 ;
  LAYER M1 ;
        RECT 15.824 6.18 15.856 6.924 ;
  LAYER M1 ;
        RECT 15.824 7.02 15.856 7.26 ;
  LAYER M1 ;
        RECT 15.824 7.356 15.856 8.1 ;
  LAYER M1 ;
        RECT 15.824 8.196 15.856 8.436 ;
  LAYER M1 ;
        RECT 15.824 8.7 15.856 8.94 ;
  LAYER M1 ;
        RECT 15.904 0.3 15.936 1.044 ;
  LAYER M1 ;
        RECT 15.904 1.476 15.936 2.22 ;
  LAYER M1 ;
        RECT 15.904 2.652 15.936 3.396 ;
  LAYER M1 ;
        RECT 15.904 3.828 15.936 4.572 ;
  LAYER M1 ;
        RECT 15.904 5.004 15.936 5.748 ;
  LAYER M1 ;
        RECT 15.904 6.18 15.936 6.924 ;
  LAYER M1 ;
        RECT 15.904 7.356 15.936 8.1 ;
  LAYER M1 ;
        RECT 15.984 0.3 16.016 1.044 ;
  LAYER M1 ;
        RECT 15.984 1.14 16.016 1.38 ;
  LAYER M1 ;
        RECT 15.984 1.476 16.016 2.22 ;
  LAYER M1 ;
        RECT 15.984 2.316 16.016 2.556 ;
  LAYER M1 ;
        RECT 15.984 2.652 16.016 3.396 ;
  LAYER M1 ;
        RECT 15.984 3.492 16.016 3.732 ;
  LAYER M1 ;
        RECT 15.984 3.828 16.016 4.572 ;
  LAYER M1 ;
        RECT 15.984 4.668 16.016 4.908 ;
  LAYER M1 ;
        RECT 15.984 5.004 16.016 5.748 ;
  LAYER M1 ;
        RECT 15.984 5.844 16.016 6.084 ;
  LAYER M1 ;
        RECT 15.984 6.18 16.016 6.924 ;
  LAYER M1 ;
        RECT 15.984 7.02 16.016 7.26 ;
  LAYER M1 ;
        RECT 15.984 7.356 16.016 8.1 ;
  LAYER M1 ;
        RECT 15.984 8.196 16.016 8.436 ;
  LAYER M1 ;
        RECT 15.984 8.7 16.016 8.94 ;
  LAYER M1 ;
        RECT 16.064 0.3 16.096 1.044 ;
  LAYER M1 ;
        RECT 16.064 1.476 16.096 2.22 ;
  LAYER M1 ;
        RECT 16.064 2.652 16.096 3.396 ;
  LAYER M1 ;
        RECT 16.064 3.828 16.096 4.572 ;
  LAYER M1 ;
        RECT 16.064 5.004 16.096 5.748 ;
  LAYER M1 ;
        RECT 16.064 6.18 16.096 6.924 ;
  LAYER M1 ;
        RECT 16.064 7.356 16.096 8.1 ;
  LAYER M2 ;
        RECT 14.124 0.32 16.116 0.352 ;
  LAYER M2 ;
        RECT 14.204 0.404 16.036 0.436 ;
  LAYER M2 ;
        RECT 14.204 1.16 16.036 1.192 ;
  LAYER M2 ;
        RECT 14.124 1.496 16.116 1.528 ;
  LAYER M2 ;
        RECT 14.204 1.58 16.036 1.612 ;
  LAYER M2 ;
        RECT 14.204 2.336 16.036 2.368 ;
  LAYER M2 ;
        RECT 14.124 2.672 16.116 2.704 ;
  LAYER M2 ;
        RECT 14.204 2.756 16.036 2.788 ;
  LAYER M2 ;
        RECT 14.204 3.512 16.036 3.544 ;
  LAYER M2 ;
        RECT 14.124 3.848 16.116 3.88 ;
  LAYER M2 ;
        RECT 14.204 3.932 16.036 3.964 ;
  LAYER M2 ;
        RECT 14.204 4.688 16.036 4.72 ;
  LAYER M2 ;
        RECT 14.124 5.024 16.116 5.056 ;
  LAYER M2 ;
        RECT 14.204 5.108 16.036 5.14 ;
  LAYER M2 ;
        RECT 14.204 5.864 16.036 5.896 ;
  LAYER M2 ;
        RECT 14.124 6.2 16.116 6.232 ;
  LAYER M2 ;
        RECT 14.204 6.284 16.036 6.316 ;
  LAYER M2 ;
        RECT 14.204 7.04 16.036 7.072 ;
  LAYER M2 ;
        RECT 14.124 7.376 16.116 7.408 ;
  LAYER M2 ;
        RECT 14.204 7.46 16.036 7.492 ;
  LAYER M2 ;
        RECT 14.204 8.216 16.036 8.248 ;
  LAYER M1 ;
        RECT 16.704 0.3 16.736 1.044 ;
  LAYER M1 ;
        RECT 16.704 1.14 16.736 1.38 ;
  LAYER M1 ;
        RECT 16.704 1.476 16.736 2.22 ;
  LAYER M1 ;
        RECT 16.704 2.316 16.736 2.556 ;
  LAYER M1 ;
        RECT 16.704 2.652 16.736 3.396 ;
  LAYER M1 ;
        RECT 16.704 3.492 16.736 3.732 ;
  LAYER M1 ;
        RECT 16.704 3.828 16.736 4.572 ;
  LAYER M1 ;
        RECT 16.704 4.668 16.736 4.908 ;
  LAYER M1 ;
        RECT 16.704 5.004 16.736 5.748 ;
  LAYER M1 ;
        RECT 16.704 5.844 16.736 6.084 ;
  LAYER M1 ;
        RECT 16.704 6.18 16.736 6.924 ;
  LAYER M1 ;
        RECT 16.704 7.02 16.736 7.26 ;
  LAYER M1 ;
        RECT 16.704 7.356 16.736 8.1 ;
  LAYER M1 ;
        RECT 16.704 8.196 16.736 8.436 ;
  LAYER M1 ;
        RECT 16.704 8.7 16.736 8.94 ;
  LAYER M1 ;
        RECT 16.624 0.3 16.656 1.044 ;
  LAYER M1 ;
        RECT 16.624 1.476 16.656 2.22 ;
  LAYER M1 ;
        RECT 16.624 2.652 16.656 3.396 ;
  LAYER M1 ;
        RECT 16.624 3.828 16.656 4.572 ;
  LAYER M1 ;
        RECT 16.624 5.004 16.656 5.748 ;
  LAYER M1 ;
        RECT 16.624 6.18 16.656 6.924 ;
  LAYER M1 ;
        RECT 16.624 7.356 16.656 8.1 ;
  LAYER M1 ;
        RECT 16.784 0.3 16.816 1.044 ;
  LAYER M1 ;
        RECT 16.784 1.476 16.816 2.22 ;
  LAYER M1 ;
        RECT 16.784 2.652 16.816 3.396 ;
  LAYER M1 ;
        RECT 16.784 3.828 16.816 4.572 ;
  LAYER M1 ;
        RECT 16.784 5.004 16.816 5.748 ;
  LAYER M1 ;
        RECT 16.784 6.18 16.816 6.924 ;
  LAYER M1 ;
        RECT 16.784 7.356 16.816 8.1 ;
  LAYER M1 ;
        RECT 16.864 0.3 16.896 1.044 ;
  LAYER M1 ;
        RECT 16.864 1.14 16.896 1.38 ;
  LAYER M1 ;
        RECT 16.864 1.476 16.896 2.22 ;
  LAYER M1 ;
        RECT 16.864 2.316 16.896 2.556 ;
  LAYER M1 ;
        RECT 16.864 2.652 16.896 3.396 ;
  LAYER M1 ;
        RECT 16.864 3.492 16.896 3.732 ;
  LAYER M1 ;
        RECT 16.864 3.828 16.896 4.572 ;
  LAYER M1 ;
        RECT 16.864 4.668 16.896 4.908 ;
  LAYER M1 ;
        RECT 16.864 5.004 16.896 5.748 ;
  LAYER M1 ;
        RECT 16.864 5.844 16.896 6.084 ;
  LAYER M1 ;
        RECT 16.864 6.18 16.896 6.924 ;
  LAYER M1 ;
        RECT 16.864 7.02 16.896 7.26 ;
  LAYER M1 ;
        RECT 16.864 7.356 16.896 8.1 ;
  LAYER M1 ;
        RECT 16.864 8.196 16.896 8.436 ;
  LAYER M1 ;
        RECT 16.864 8.7 16.896 8.94 ;
  LAYER M1 ;
        RECT 16.944 0.3 16.976 1.044 ;
  LAYER M1 ;
        RECT 16.944 1.476 16.976 2.22 ;
  LAYER M1 ;
        RECT 16.944 2.652 16.976 3.396 ;
  LAYER M1 ;
        RECT 16.944 3.828 16.976 4.572 ;
  LAYER M1 ;
        RECT 16.944 5.004 16.976 5.748 ;
  LAYER M1 ;
        RECT 16.944 6.18 16.976 6.924 ;
  LAYER M1 ;
        RECT 16.944 7.356 16.976 8.1 ;
  LAYER M1 ;
        RECT 17.024 0.3 17.056 1.044 ;
  LAYER M1 ;
        RECT 17.024 1.14 17.056 1.38 ;
  LAYER M1 ;
        RECT 17.024 1.476 17.056 2.22 ;
  LAYER M1 ;
        RECT 17.024 2.316 17.056 2.556 ;
  LAYER M1 ;
        RECT 17.024 2.652 17.056 3.396 ;
  LAYER M1 ;
        RECT 17.024 3.492 17.056 3.732 ;
  LAYER M1 ;
        RECT 17.024 3.828 17.056 4.572 ;
  LAYER M1 ;
        RECT 17.024 4.668 17.056 4.908 ;
  LAYER M1 ;
        RECT 17.024 5.004 17.056 5.748 ;
  LAYER M1 ;
        RECT 17.024 5.844 17.056 6.084 ;
  LAYER M1 ;
        RECT 17.024 6.18 17.056 6.924 ;
  LAYER M1 ;
        RECT 17.024 7.02 17.056 7.26 ;
  LAYER M1 ;
        RECT 17.024 7.356 17.056 8.1 ;
  LAYER M1 ;
        RECT 17.024 8.196 17.056 8.436 ;
  LAYER M1 ;
        RECT 17.024 8.7 17.056 8.94 ;
  LAYER M1 ;
        RECT 17.104 0.3 17.136 1.044 ;
  LAYER M1 ;
        RECT 17.104 1.476 17.136 2.22 ;
  LAYER M1 ;
        RECT 17.104 2.652 17.136 3.396 ;
  LAYER M1 ;
        RECT 17.104 3.828 17.136 4.572 ;
  LAYER M1 ;
        RECT 17.104 5.004 17.136 5.748 ;
  LAYER M1 ;
        RECT 17.104 6.18 17.136 6.924 ;
  LAYER M1 ;
        RECT 17.104 7.356 17.136 8.1 ;
  LAYER M1 ;
        RECT 17.184 0.3 17.216 1.044 ;
  LAYER M1 ;
        RECT 17.184 1.14 17.216 1.38 ;
  LAYER M1 ;
        RECT 17.184 1.476 17.216 2.22 ;
  LAYER M1 ;
        RECT 17.184 2.316 17.216 2.556 ;
  LAYER M1 ;
        RECT 17.184 2.652 17.216 3.396 ;
  LAYER M1 ;
        RECT 17.184 3.492 17.216 3.732 ;
  LAYER M1 ;
        RECT 17.184 3.828 17.216 4.572 ;
  LAYER M1 ;
        RECT 17.184 4.668 17.216 4.908 ;
  LAYER M1 ;
        RECT 17.184 5.004 17.216 5.748 ;
  LAYER M1 ;
        RECT 17.184 5.844 17.216 6.084 ;
  LAYER M1 ;
        RECT 17.184 6.18 17.216 6.924 ;
  LAYER M1 ;
        RECT 17.184 7.02 17.216 7.26 ;
  LAYER M1 ;
        RECT 17.184 7.356 17.216 8.1 ;
  LAYER M1 ;
        RECT 17.184 8.196 17.216 8.436 ;
  LAYER M1 ;
        RECT 17.184 8.7 17.216 8.94 ;
  LAYER M1 ;
        RECT 17.264 0.3 17.296 1.044 ;
  LAYER M1 ;
        RECT 17.264 1.476 17.296 2.22 ;
  LAYER M1 ;
        RECT 17.264 2.652 17.296 3.396 ;
  LAYER M1 ;
        RECT 17.264 3.828 17.296 4.572 ;
  LAYER M1 ;
        RECT 17.264 5.004 17.296 5.748 ;
  LAYER M1 ;
        RECT 17.264 6.18 17.296 6.924 ;
  LAYER M1 ;
        RECT 17.264 7.356 17.296 8.1 ;
  LAYER M1 ;
        RECT 17.344 0.3 17.376 1.044 ;
  LAYER M1 ;
        RECT 17.344 1.14 17.376 1.38 ;
  LAYER M1 ;
        RECT 17.344 1.476 17.376 2.22 ;
  LAYER M1 ;
        RECT 17.344 2.316 17.376 2.556 ;
  LAYER M1 ;
        RECT 17.344 2.652 17.376 3.396 ;
  LAYER M1 ;
        RECT 17.344 3.492 17.376 3.732 ;
  LAYER M1 ;
        RECT 17.344 3.828 17.376 4.572 ;
  LAYER M1 ;
        RECT 17.344 4.668 17.376 4.908 ;
  LAYER M1 ;
        RECT 17.344 5.004 17.376 5.748 ;
  LAYER M1 ;
        RECT 17.344 5.844 17.376 6.084 ;
  LAYER M1 ;
        RECT 17.344 6.18 17.376 6.924 ;
  LAYER M1 ;
        RECT 17.344 7.02 17.376 7.26 ;
  LAYER M1 ;
        RECT 17.344 7.356 17.376 8.1 ;
  LAYER M1 ;
        RECT 17.344 8.196 17.376 8.436 ;
  LAYER M1 ;
        RECT 17.344 8.7 17.376 8.94 ;
  LAYER M1 ;
        RECT 17.424 0.3 17.456 1.044 ;
  LAYER M1 ;
        RECT 17.424 1.476 17.456 2.22 ;
  LAYER M1 ;
        RECT 17.424 2.652 17.456 3.396 ;
  LAYER M1 ;
        RECT 17.424 3.828 17.456 4.572 ;
  LAYER M1 ;
        RECT 17.424 5.004 17.456 5.748 ;
  LAYER M1 ;
        RECT 17.424 6.18 17.456 6.924 ;
  LAYER M1 ;
        RECT 17.424 7.356 17.456 8.1 ;
  LAYER M1 ;
        RECT 17.504 0.3 17.536 1.044 ;
  LAYER M1 ;
        RECT 17.504 1.14 17.536 1.38 ;
  LAYER M1 ;
        RECT 17.504 1.476 17.536 2.22 ;
  LAYER M1 ;
        RECT 17.504 2.316 17.536 2.556 ;
  LAYER M1 ;
        RECT 17.504 2.652 17.536 3.396 ;
  LAYER M1 ;
        RECT 17.504 3.492 17.536 3.732 ;
  LAYER M1 ;
        RECT 17.504 3.828 17.536 4.572 ;
  LAYER M1 ;
        RECT 17.504 4.668 17.536 4.908 ;
  LAYER M1 ;
        RECT 17.504 5.004 17.536 5.748 ;
  LAYER M1 ;
        RECT 17.504 5.844 17.536 6.084 ;
  LAYER M1 ;
        RECT 17.504 6.18 17.536 6.924 ;
  LAYER M1 ;
        RECT 17.504 7.02 17.536 7.26 ;
  LAYER M1 ;
        RECT 17.504 7.356 17.536 8.1 ;
  LAYER M1 ;
        RECT 17.504 8.196 17.536 8.436 ;
  LAYER M1 ;
        RECT 17.504 8.7 17.536 8.94 ;
  LAYER M1 ;
        RECT 17.584 0.3 17.616 1.044 ;
  LAYER M1 ;
        RECT 17.584 1.476 17.616 2.22 ;
  LAYER M1 ;
        RECT 17.584 2.652 17.616 3.396 ;
  LAYER M1 ;
        RECT 17.584 3.828 17.616 4.572 ;
  LAYER M1 ;
        RECT 17.584 5.004 17.616 5.748 ;
  LAYER M1 ;
        RECT 17.584 6.18 17.616 6.924 ;
  LAYER M1 ;
        RECT 17.584 7.356 17.616 8.1 ;
  LAYER M1 ;
        RECT 17.664 0.3 17.696 1.044 ;
  LAYER M1 ;
        RECT 17.664 1.14 17.696 1.38 ;
  LAYER M1 ;
        RECT 17.664 1.476 17.696 2.22 ;
  LAYER M1 ;
        RECT 17.664 2.316 17.696 2.556 ;
  LAYER M1 ;
        RECT 17.664 2.652 17.696 3.396 ;
  LAYER M1 ;
        RECT 17.664 3.492 17.696 3.732 ;
  LAYER M1 ;
        RECT 17.664 3.828 17.696 4.572 ;
  LAYER M1 ;
        RECT 17.664 4.668 17.696 4.908 ;
  LAYER M1 ;
        RECT 17.664 5.004 17.696 5.748 ;
  LAYER M1 ;
        RECT 17.664 5.844 17.696 6.084 ;
  LAYER M1 ;
        RECT 17.664 6.18 17.696 6.924 ;
  LAYER M1 ;
        RECT 17.664 7.02 17.696 7.26 ;
  LAYER M1 ;
        RECT 17.664 7.356 17.696 8.1 ;
  LAYER M1 ;
        RECT 17.664 8.196 17.696 8.436 ;
  LAYER M1 ;
        RECT 17.664 8.7 17.696 8.94 ;
  LAYER M1 ;
        RECT 17.744 0.3 17.776 1.044 ;
  LAYER M1 ;
        RECT 17.744 1.476 17.776 2.22 ;
  LAYER M1 ;
        RECT 17.744 2.652 17.776 3.396 ;
  LAYER M1 ;
        RECT 17.744 3.828 17.776 4.572 ;
  LAYER M1 ;
        RECT 17.744 5.004 17.776 5.748 ;
  LAYER M1 ;
        RECT 17.744 6.18 17.776 6.924 ;
  LAYER M1 ;
        RECT 17.744 7.356 17.776 8.1 ;
  LAYER M1 ;
        RECT 17.824 0.3 17.856 1.044 ;
  LAYER M1 ;
        RECT 17.824 1.14 17.856 1.38 ;
  LAYER M1 ;
        RECT 17.824 1.476 17.856 2.22 ;
  LAYER M1 ;
        RECT 17.824 2.316 17.856 2.556 ;
  LAYER M1 ;
        RECT 17.824 2.652 17.856 3.396 ;
  LAYER M1 ;
        RECT 17.824 3.492 17.856 3.732 ;
  LAYER M1 ;
        RECT 17.824 3.828 17.856 4.572 ;
  LAYER M1 ;
        RECT 17.824 4.668 17.856 4.908 ;
  LAYER M1 ;
        RECT 17.824 5.004 17.856 5.748 ;
  LAYER M1 ;
        RECT 17.824 5.844 17.856 6.084 ;
  LAYER M1 ;
        RECT 17.824 6.18 17.856 6.924 ;
  LAYER M1 ;
        RECT 17.824 7.02 17.856 7.26 ;
  LAYER M1 ;
        RECT 17.824 7.356 17.856 8.1 ;
  LAYER M1 ;
        RECT 17.824 8.196 17.856 8.436 ;
  LAYER M1 ;
        RECT 17.824 8.7 17.856 8.94 ;
  LAYER M1 ;
        RECT 17.904 0.3 17.936 1.044 ;
  LAYER M1 ;
        RECT 17.904 1.476 17.936 2.22 ;
  LAYER M1 ;
        RECT 17.904 2.652 17.936 3.396 ;
  LAYER M1 ;
        RECT 17.904 3.828 17.936 4.572 ;
  LAYER M1 ;
        RECT 17.904 5.004 17.936 5.748 ;
  LAYER M1 ;
        RECT 17.904 6.18 17.936 6.924 ;
  LAYER M1 ;
        RECT 17.904 7.356 17.936 8.1 ;
  LAYER M1 ;
        RECT 17.984 0.3 18.016 1.044 ;
  LAYER M1 ;
        RECT 17.984 1.14 18.016 1.38 ;
  LAYER M1 ;
        RECT 17.984 1.476 18.016 2.22 ;
  LAYER M1 ;
        RECT 17.984 2.316 18.016 2.556 ;
  LAYER M1 ;
        RECT 17.984 2.652 18.016 3.396 ;
  LAYER M1 ;
        RECT 17.984 3.492 18.016 3.732 ;
  LAYER M1 ;
        RECT 17.984 3.828 18.016 4.572 ;
  LAYER M1 ;
        RECT 17.984 4.668 18.016 4.908 ;
  LAYER M1 ;
        RECT 17.984 5.004 18.016 5.748 ;
  LAYER M1 ;
        RECT 17.984 5.844 18.016 6.084 ;
  LAYER M1 ;
        RECT 17.984 6.18 18.016 6.924 ;
  LAYER M1 ;
        RECT 17.984 7.02 18.016 7.26 ;
  LAYER M1 ;
        RECT 17.984 7.356 18.016 8.1 ;
  LAYER M1 ;
        RECT 17.984 8.196 18.016 8.436 ;
  LAYER M1 ;
        RECT 17.984 8.7 18.016 8.94 ;
  LAYER M1 ;
        RECT 18.064 0.3 18.096 1.044 ;
  LAYER M1 ;
        RECT 18.064 1.476 18.096 2.22 ;
  LAYER M1 ;
        RECT 18.064 2.652 18.096 3.396 ;
  LAYER M1 ;
        RECT 18.064 3.828 18.096 4.572 ;
  LAYER M1 ;
        RECT 18.064 5.004 18.096 5.748 ;
  LAYER M1 ;
        RECT 18.064 6.18 18.096 6.924 ;
  LAYER M1 ;
        RECT 18.064 7.356 18.096 8.1 ;
  LAYER M1 ;
        RECT 18.144 0.3 18.176 1.044 ;
  LAYER M1 ;
        RECT 18.144 1.14 18.176 1.38 ;
  LAYER M1 ;
        RECT 18.144 1.476 18.176 2.22 ;
  LAYER M1 ;
        RECT 18.144 2.316 18.176 2.556 ;
  LAYER M1 ;
        RECT 18.144 2.652 18.176 3.396 ;
  LAYER M1 ;
        RECT 18.144 3.492 18.176 3.732 ;
  LAYER M1 ;
        RECT 18.144 3.828 18.176 4.572 ;
  LAYER M1 ;
        RECT 18.144 4.668 18.176 4.908 ;
  LAYER M1 ;
        RECT 18.144 5.004 18.176 5.748 ;
  LAYER M1 ;
        RECT 18.144 5.844 18.176 6.084 ;
  LAYER M1 ;
        RECT 18.144 6.18 18.176 6.924 ;
  LAYER M1 ;
        RECT 18.144 7.02 18.176 7.26 ;
  LAYER M1 ;
        RECT 18.144 7.356 18.176 8.1 ;
  LAYER M1 ;
        RECT 18.144 8.196 18.176 8.436 ;
  LAYER M1 ;
        RECT 18.144 8.7 18.176 8.94 ;
  LAYER M1 ;
        RECT 18.224 0.3 18.256 1.044 ;
  LAYER M1 ;
        RECT 18.224 1.476 18.256 2.22 ;
  LAYER M1 ;
        RECT 18.224 2.652 18.256 3.396 ;
  LAYER M1 ;
        RECT 18.224 3.828 18.256 4.572 ;
  LAYER M1 ;
        RECT 18.224 5.004 18.256 5.748 ;
  LAYER M1 ;
        RECT 18.224 6.18 18.256 6.924 ;
  LAYER M1 ;
        RECT 18.224 7.356 18.256 8.1 ;
  LAYER M1 ;
        RECT 18.304 0.3 18.336 1.044 ;
  LAYER M1 ;
        RECT 18.304 1.14 18.336 1.38 ;
  LAYER M1 ;
        RECT 18.304 1.476 18.336 2.22 ;
  LAYER M1 ;
        RECT 18.304 2.316 18.336 2.556 ;
  LAYER M1 ;
        RECT 18.304 2.652 18.336 3.396 ;
  LAYER M1 ;
        RECT 18.304 3.492 18.336 3.732 ;
  LAYER M1 ;
        RECT 18.304 3.828 18.336 4.572 ;
  LAYER M1 ;
        RECT 18.304 4.668 18.336 4.908 ;
  LAYER M1 ;
        RECT 18.304 5.004 18.336 5.748 ;
  LAYER M1 ;
        RECT 18.304 5.844 18.336 6.084 ;
  LAYER M1 ;
        RECT 18.304 6.18 18.336 6.924 ;
  LAYER M1 ;
        RECT 18.304 7.02 18.336 7.26 ;
  LAYER M1 ;
        RECT 18.304 7.356 18.336 8.1 ;
  LAYER M1 ;
        RECT 18.304 8.196 18.336 8.436 ;
  LAYER M1 ;
        RECT 18.304 8.7 18.336 8.94 ;
  LAYER M1 ;
        RECT 18.384 0.3 18.416 1.044 ;
  LAYER M1 ;
        RECT 18.384 1.476 18.416 2.22 ;
  LAYER M1 ;
        RECT 18.384 2.652 18.416 3.396 ;
  LAYER M1 ;
        RECT 18.384 3.828 18.416 4.572 ;
  LAYER M1 ;
        RECT 18.384 5.004 18.416 5.748 ;
  LAYER M1 ;
        RECT 18.384 6.18 18.416 6.924 ;
  LAYER M1 ;
        RECT 18.384 7.356 18.416 8.1 ;
  LAYER M1 ;
        RECT 18.464 0.3 18.496 1.044 ;
  LAYER M1 ;
        RECT 18.464 1.14 18.496 1.38 ;
  LAYER M1 ;
        RECT 18.464 1.476 18.496 2.22 ;
  LAYER M1 ;
        RECT 18.464 2.316 18.496 2.556 ;
  LAYER M1 ;
        RECT 18.464 2.652 18.496 3.396 ;
  LAYER M1 ;
        RECT 18.464 3.492 18.496 3.732 ;
  LAYER M1 ;
        RECT 18.464 3.828 18.496 4.572 ;
  LAYER M1 ;
        RECT 18.464 4.668 18.496 4.908 ;
  LAYER M1 ;
        RECT 18.464 5.004 18.496 5.748 ;
  LAYER M1 ;
        RECT 18.464 5.844 18.496 6.084 ;
  LAYER M1 ;
        RECT 18.464 6.18 18.496 6.924 ;
  LAYER M1 ;
        RECT 18.464 7.02 18.496 7.26 ;
  LAYER M1 ;
        RECT 18.464 7.356 18.496 8.1 ;
  LAYER M1 ;
        RECT 18.464 8.196 18.496 8.436 ;
  LAYER M1 ;
        RECT 18.464 8.7 18.496 8.94 ;
  LAYER M1 ;
        RECT 18.544 0.3 18.576 1.044 ;
  LAYER M1 ;
        RECT 18.544 1.476 18.576 2.22 ;
  LAYER M1 ;
        RECT 18.544 2.652 18.576 3.396 ;
  LAYER M1 ;
        RECT 18.544 3.828 18.576 4.572 ;
  LAYER M1 ;
        RECT 18.544 5.004 18.576 5.748 ;
  LAYER M1 ;
        RECT 18.544 6.18 18.576 6.924 ;
  LAYER M1 ;
        RECT 18.544 7.356 18.576 8.1 ;
  LAYER M1 ;
        RECT 18.624 0.3 18.656 1.044 ;
  LAYER M1 ;
        RECT 18.624 1.14 18.656 1.38 ;
  LAYER M1 ;
        RECT 18.624 1.476 18.656 2.22 ;
  LAYER M1 ;
        RECT 18.624 2.316 18.656 2.556 ;
  LAYER M1 ;
        RECT 18.624 2.652 18.656 3.396 ;
  LAYER M1 ;
        RECT 18.624 3.492 18.656 3.732 ;
  LAYER M1 ;
        RECT 18.624 3.828 18.656 4.572 ;
  LAYER M1 ;
        RECT 18.624 4.668 18.656 4.908 ;
  LAYER M1 ;
        RECT 18.624 5.004 18.656 5.748 ;
  LAYER M1 ;
        RECT 18.624 5.844 18.656 6.084 ;
  LAYER M1 ;
        RECT 18.624 6.18 18.656 6.924 ;
  LAYER M1 ;
        RECT 18.624 7.02 18.656 7.26 ;
  LAYER M1 ;
        RECT 18.624 7.356 18.656 8.1 ;
  LAYER M1 ;
        RECT 18.624 8.196 18.656 8.436 ;
  LAYER M1 ;
        RECT 18.624 8.7 18.656 8.94 ;
  LAYER M1 ;
        RECT 18.704 0.3 18.736 1.044 ;
  LAYER M1 ;
        RECT 18.704 1.476 18.736 2.22 ;
  LAYER M1 ;
        RECT 18.704 2.652 18.736 3.396 ;
  LAYER M1 ;
        RECT 18.704 3.828 18.736 4.572 ;
  LAYER M1 ;
        RECT 18.704 5.004 18.736 5.748 ;
  LAYER M1 ;
        RECT 18.704 6.18 18.736 6.924 ;
  LAYER M1 ;
        RECT 18.704 7.356 18.736 8.1 ;
  LAYER M1 ;
        RECT 18.784 0.3 18.816 1.044 ;
  LAYER M1 ;
        RECT 18.784 1.14 18.816 1.38 ;
  LAYER M1 ;
        RECT 18.784 1.476 18.816 2.22 ;
  LAYER M1 ;
        RECT 18.784 2.316 18.816 2.556 ;
  LAYER M1 ;
        RECT 18.784 2.652 18.816 3.396 ;
  LAYER M1 ;
        RECT 18.784 3.492 18.816 3.732 ;
  LAYER M1 ;
        RECT 18.784 3.828 18.816 4.572 ;
  LAYER M1 ;
        RECT 18.784 4.668 18.816 4.908 ;
  LAYER M1 ;
        RECT 18.784 5.004 18.816 5.748 ;
  LAYER M1 ;
        RECT 18.784 5.844 18.816 6.084 ;
  LAYER M1 ;
        RECT 18.784 6.18 18.816 6.924 ;
  LAYER M1 ;
        RECT 18.784 7.02 18.816 7.26 ;
  LAYER M1 ;
        RECT 18.784 7.356 18.816 8.1 ;
  LAYER M1 ;
        RECT 18.784 8.196 18.816 8.436 ;
  LAYER M1 ;
        RECT 18.784 8.7 18.816 8.94 ;
  LAYER M1 ;
        RECT 18.864 0.3 18.896 1.044 ;
  LAYER M1 ;
        RECT 18.864 1.476 18.896 2.22 ;
  LAYER M1 ;
        RECT 18.864 2.652 18.896 3.396 ;
  LAYER M1 ;
        RECT 18.864 3.828 18.896 4.572 ;
  LAYER M1 ;
        RECT 18.864 5.004 18.896 5.748 ;
  LAYER M1 ;
        RECT 18.864 6.18 18.896 6.924 ;
  LAYER M1 ;
        RECT 18.864 7.356 18.896 8.1 ;
  LAYER M1 ;
        RECT 18.944 0.3 18.976 1.044 ;
  LAYER M1 ;
        RECT 18.944 1.14 18.976 1.38 ;
  LAYER M1 ;
        RECT 18.944 1.476 18.976 2.22 ;
  LAYER M1 ;
        RECT 18.944 2.316 18.976 2.556 ;
  LAYER M1 ;
        RECT 18.944 2.652 18.976 3.396 ;
  LAYER M1 ;
        RECT 18.944 3.492 18.976 3.732 ;
  LAYER M1 ;
        RECT 18.944 3.828 18.976 4.572 ;
  LAYER M1 ;
        RECT 18.944 4.668 18.976 4.908 ;
  LAYER M1 ;
        RECT 18.944 5.004 18.976 5.748 ;
  LAYER M1 ;
        RECT 18.944 5.844 18.976 6.084 ;
  LAYER M1 ;
        RECT 18.944 6.18 18.976 6.924 ;
  LAYER M1 ;
        RECT 18.944 7.02 18.976 7.26 ;
  LAYER M1 ;
        RECT 18.944 7.356 18.976 8.1 ;
  LAYER M1 ;
        RECT 18.944 8.196 18.976 8.436 ;
  LAYER M1 ;
        RECT 18.944 8.7 18.976 8.94 ;
  LAYER M1 ;
        RECT 19.024 0.3 19.056 1.044 ;
  LAYER M1 ;
        RECT 19.024 1.476 19.056 2.22 ;
  LAYER M1 ;
        RECT 19.024 2.652 19.056 3.396 ;
  LAYER M1 ;
        RECT 19.024 3.828 19.056 4.572 ;
  LAYER M1 ;
        RECT 19.024 5.004 19.056 5.748 ;
  LAYER M1 ;
        RECT 19.024 6.18 19.056 6.924 ;
  LAYER M1 ;
        RECT 19.024 7.356 19.056 8.1 ;
  LAYER M1 ;
        RECT 19.104 0.3 19.136 1.044 ;
  LAYER M1 ;
        RECT 19.104 1.14 19.136 1.38 ;
  LAYER M1 ;
        RECT 19.104 1.476 19.136 2.22 ;
  LAYER M1 ;
        RECT 19.104 2.316 19.136 2.556 ;
  LAYER M1 ;
        RECT 19.104 2.652 19.136 3.396 ;
  LAYER M1 ;
        RECT 19.104 3.492 19.136 3.732 ;
  LAYER M1 ;
        RECT 19.104 3.828 19.136 4.572 ;
  LAYER M1 ;
        RECT 19.104 4.668 19.136 4.908 ;
  LAYER M1 ;
        RECT 19.104 5.004 19.136 5.748 ;
  LAYER M1 ;
        RECT 19.104 5.844 19.136 6.084 ;
  LAYER M1 ;
        RECT 19.104 6.18 19.136 6.924 ;
  LAYER M1 ;
        RECT 19.104 7.02 19.136 7.26 ;
  LAYER M1 ;
        RECT 19.104 7.356 19.136 8.1 ;
  LAYER M1 ;
        RECT 19.104 8.196 19.136 8.436 ;
  LAYER M1 ;
        RECT 19.104 8.7 19.136 8.94 ;
  LAYER M1 ;
        RECT 19.184 0.3 19.216 1.044 ;
  LAYER M1 ;
        RECT 19.184 1.476 19.216 2.22 ;
  LAYER M1 ;
        RECT 19.184 2.652 19.216 3.396 ;
  LAYER M1 ;
        RECT 19.184 3.828 19.216 4.572 ;
  LAYER M1 ;
        RECT 19.184 5.004 19.216 5.748 ;
  LAYER M1 ;
        RECT 19.184 6.18 19.216 6.924 ;
  LAYER M1 ;
        RECT 19.184 7.356 19.216 8.1 ;
  LAYER M1 ;
        RECT 19.264 0.3 19.296 1.044 ;
  LAYER M1 ;
        RECT 19.264 1.14 19.296 1.38 ;
  LAYER M1 ;
        RECT 19.264 1.476 19.296 2.22 ;
  LAYER M1 ;
        RECT 19.264 2.316 19.296 2.556 ;
  LAYER M1 ;
        RECT 19.264 2.652 19.296 3.396 ;
  LAYER M1 ;
        RECT 19.264 3.492 19.296 3.732 ;
  LAYER M1 ;
        RECT 19.264 3.828 19.296 4.572 ;
  LAYER M1 ;
        RECT 19.264 4.668 19.296 4.908 ;
  LAYER M1 ;
        RECT 19.264 5.004 19.296 5.748 ;
  LAYER M1 ;
        RECT 19.264 5.844 19.296 6.084 ;
  LAYER M1 ;
        RECT 19.264 6.18 19.296 6.924 ;
  LAYER M1 ;
        RECT 19.264 7.02 19.296 7.26 ;
  LAYER M1 ;
        RECT 19.264 7.356 19.296 8.1 ;
  LAYER M1 ;
        RECT 19.264 8.196 19.296 8.436 ;
  LAYER M1 ;
        RECT 19.264 8.7 19.296 8.94 ;
  LAYER M1 ;
        RECT 19.344 0.3 19.376 1.044 ;
  LAYER M1 ;
        RECT 19.344 1.476 19.376 2.22 ;
  LAYER M1 ;
        RECT 19.344 2.652 19.376 3.396 ;
  LAYER M1 ;
        RECT 19.344 3.828 19.376 4.572 ;
  LAYER M1 ;
        RECT 19.344 5.004 19.376 5.748 ;
  LAYER M1 ;
        RECT 19.344 6.18 19.376 6.924 ;
  LAYER M1 ;
        RECT 19.344 7.356 19.376 8.1 ;
  LAYER M1 ;
        RECT 19.424 0.3 19.456 1.044 ;
  LAYER M1 ;
        RECT 19.424 1.14 19.456 1.38 ;
  LAYER M1 ;
        RECT 19.424 1.476 19.456 2.22 ;
  LAYER M1 ;
        RECT 19.424 2.316 19.456 2.556 ;
  LAYER M1 ;
        RECT 19.424 2.652 19.456 3.396 ;
  LAYER M1 ;
        RECT 19.424 3.492 19.456 3.732 ;
  LAYER M1 ;
        RECT 19.424 3.828 19.456 4.572 ;
  LAYER M1 ;
        RECT 19.424 4.668 19.456 4.908 ;
  LAYER M1 ;
        RECT 19.424 5.004 19.456 5.748 ;
  LAYER M1 ;
        RECT 19.424 5.844 19.456 6.084 ;
  LAYER M1 ;
        RECT 19.424 6.18 19.456 6.924 ;
  LAYER M1 ;
        RECT 19.424 7.02 19.456 7.26 ;
  LAYER M1 ;
        RECT 19.424 7.356 19.456 8.1 ;
  LAYER M1 ;
        RECT 19.424 8.196 19.456 8.436 ;
  LAYER M1 ;
        RECT 19.424 8.7 19.456 8.94 ;
  LAYER M1 ;
        RECT 19.504 0.3 19.536 1.044 ;
  LAYER M1 ;
        RECT 19.504 1.476 19.536 2.22 ;
  LAYER M1 ;
        RECT 19.504 2.652 19.536 3.396 ;
  LAYER M1 ;
        RECT 19.504 3.828 19.536 4.572 ;
  LAYER M1 ;
        RECT 19.504 5.004 19.536 5.748 ;
  LAYER M1 ;
        RECT 19.504 6.18 19.536 6.924 ;
  LAYER M1 ;
        RECT 19.504 7.356 19.536 8.1 ;
  LAYER M1 ;
        RECT 19.584 0.3 19.616 1.044 ;
  LAYER M1 ;
        RECT 19.584 1.14 19.616 1.38 ;
  LAYER M1 ;
        RECT 19.584 1.476 19.616 2.22 ;
  LAYER M1 ;
        RECT 19.584 2.316 19.616 2.556 ;
  LAYER M1 ;
        RECT 19.584 2.652 19.616 3.396 ;
  LAYER M1 ;
        RECT 19.584 3.492 19.616 3.732 ;
  LAYER M1 ;
        RECT 19.584 3.828 19.616 4.572 ;
  LAYER M1 ;
        RECT 19.584 4.668 19.616 4.908 ;
  LAYER M1 ;
        RECT 19.584 5.004 19.616 5.748 ;
  LAYER M1 ;
        RECT 19.584 5.844 19.616 6.084 ;
  LAYER M1 ;
        RECT 19.584 6.18 19.616 6.924 ;
  LAYER M1 ;
        RECT 19.584 7.02 19.616 7.26 ;
  LAYER M1 ;
        RECT 19.584 7.356 19.616 8.1 ;
  LAYER M1 ;
        RECT 19.584 8.196 19.616 8.436 ;
  LAYER M1 ;
        RECT 19.584 8.7 19.616 8.94 ;
  LAYER M1 ;
        RECT 19.664 0.3 19.696 1.044 ;
  LAYER M1 ;
        RECT 19.664 1.476 19.696 2.22 ;
  LAYER M1 ;
        RECT 19.664 2.652 19.696 3.396 ;
  LAYER M1 ;
        RECT 19.664 3.828 19.696 4.572 ;
  LAYER M1 ;
        RECT 19.664 5.004 19.696 5.748 ;
  LAYER M1 ;
        RECT 19.664 6.18 19.696 6.924 ;
  LAYER M1 ;
        RECT 19.664 7.356 19.696 8.1 ;
  LAYER M1 ;
        RECT 19.744 0.3 19.776 1.044 ;
  LAYER M1 ;
        RECT 19.744 1.14 19.776 1.38 ;
  LAYER M1 ;
        RECT 19.744 1.476 19.776 2.22 ;
  LAYER M1 ;
        RECT 19.744 2.316 19.776 2.556 ;
  LAYER M1 ;
        RECT 19.744 2.652 19.776 3.396 ;
  LAYER M1 ;
        RECT 19.744 3.492 19.776 3.732 ;
  LAYER M1 ;
        RECT 19.744 3.828 19.776 4.572 ;
  LAYER M1 ;
        RECT 19.744 4.668 19.776 4.908 ;
  LAYER M1 ;
        RECT 19.744 5.004 19.776 5.748 ;
  LAYER M1 ;
        RECT 19.744 5.844 19.776 6.084 ;
  LAYER M1 ;
        RECT 19.744 6.18 19.776 6.924 ;
  LAYER M1 ;
        RECT 19.744 7.02 19.776 7.26 ;
  LAYER M1 ;
        RECT 19.744 7.356 19.776 8.1 ;
  LAYER M1 ;
        RECT 19.744 8.196 19.776 8.436 ;
  LAYER M1 ;
        RECT 19.744 8.7 19.776 8.94 ;
  LAYER M1 ;
        RECT 19.824 0.3 19.856 1.044 ;
  LAYER M1 ;
        RECT 19.824 1.476 19.856 2.22 ;
  LAYER M1 ;
        RECT 19.824 2.652 19.856 3.396 ;
  LAYER M1 ;
        RECT 19.824 3.828 19.856 4.572 ;
  LAYER M1 ;
        RECT 19.824 5.004 19.856 5.748 ;
  LAYER M1 ;
        RECT 19.824 6.18 19.856 6.924 ;
  LAYER M1 ;
        RECT 19.824 7.356 19.856 8.1 ;
  LAYER M1 ;
        RECT 19.904 0.3 19.936 1.044 ;
  LAYER M1 ;
        RECT 19.904 1.14 19.936 1.38 ;
  LAYER M1 ;
        RECT 19.904 1.476 19.936 2.22 ;
  LAYER M1 ;
        RECT 19.904 2.316 19.936 2.556 ;
  LAYER M1 ;
        RECT 19.904 2.652 19.936 3.396 ;
  LAYER M1 ;
        RECT 19.904 3.492 19.936 3.732 ;
  LAYER M1 ;
        RECT 19.904 3.828 19.936 4.572 ;
  LAYER M1 ;
        RECT 19.904 4.668 19.936 4.908 ;
  LAYER M1 ;
        RECT 19.904 5.004 19.936 5.748 ;
  LAYER M1 ;
        RECT 19.904 5.844 19.936 6.084 ;
  LAYER M1 ;
        RECT 19.904 6.18 19.936 6.924 ;
  LAYER M1 ;
        RECT 19.904 7.02 19.936 7.26 ;
  LAYER M1 ;
        RECT 19.904 7.356 19.936 8.1 ;
  LAYER M1 ;
        RECT 19.904 8.196 19.936 8.436 ;
  LAYER M1 ;
        RECT 19.904 8.7 19.936 8.94 ;
  LAYER M1 ;
        RECT 19.984 0.3 20.016 1.044 ;
  LAYER M1 ;
        RECT 19.984 1.476 20.016 2.22 ;
  LAYER M1 ;
        RECT 19.984 2.652 20.016 3.396 ;
  LAYER M1 ;
        RECT 19.984 3.828 20.016 4.572 ;
  LAYER M1 ;
        RECT 19.984 5.004 20.016 5.748 ;
  LAYER M1 ;
        RECT 19.984 6.18 20.016 6.924 ;
  LAYER M1 ;
        RECT 19.984 7.356 20.016 8.1 ;
  LAYER M1 ;
        RECT 20.064 0.3 20.096 1.044 ;
  LAYER M1 ;
        RECT 20.064 1.14 20.096 1.38 ;
  LAYER M1 ;
        RECT 20.064 1.476 20.096 2.22 ;
  LAYER M1 ;
        RECT 20.064 2.316 20.096 2.556 ;
  LAYER M1 ;
        RECT 20.064 2.652 20.096 3.396 ;
  LAYER M1 ;
        RECT 20.064 3.492 20.096 3.732 ;
  LAYER M1 ;
        RECT 20.064 3.828 20.096 4.572 ;
  LAYER M1 ;
        RECT 20.064 4.668 20.096 4.908 ;
  LAYER M1 ;
        RECT 20.064 5.004 20.096 5.748 ;
  LAYER M1 ;
        RECT 20.064 5.844 20.096 6.084 ;
  LAYER M1 ;
        RECT 20.064 6.18 20.096 6.924 ;
  LAYER M1 ;
        RECT 20.064 7.02 20.096 7.26 ;
  LAYER M1 ;
        RECT 20.064 7.356 20.096 8.1 ;
  LAYER M1 ;
        RECT 20.064 8.196 20.096 8.436 ;
  LAYER M1 ;
        RECT 20.064 8.7 20.096 8.94 ;
  LAYER M1 ;
        RECT 20.144 0.3 20.176 1.044 ;
  LAYER M1 ;
        RECT 20.144 1.476 20.176 2.22 ;
  LAYER M1 ;
        RECT 20.144 2.652 20.176 3.396 ;
  LAYER M1 ;
        RECT 20.144 3.828 20.176 4.572 ;
  LAYER M1 ;
        RECT 20.144 5.004 20.176 5.748 ;
  LAYER M1 ;
        RECT 20.144 6.18 20.176 6.924 ;
  LAYER M1 ;
        RECT 20.144 7.356 20.176 8.1 ;
  LAYER M1 ;
        RECT 20.224 0.3 20.256 1.044 ;
  LAYER M1 ;
        RECT 20.224 1.14 20.256 1.38 ;
  LAYER M1 ;
        RECT 20.224 1.476 20.256 2.22 ;
  LAYER M1 ;
        RECT 20.224 2.316 20.256 2.556 ;
  LAYER M1 ;
        RECT 20.224 2.652 20.256 3.396 ;
  LAYER M1 ;
        RECT 20.224 3.492 20.256 3.732 ;
  LAYER M1 ;
        RECT 20.224 3.828 20.256 4.572 ;
  LAYER M1 ;
        RECT 20.224 4.668 20.256 4.908 ;
  LAYER M1 ;
        RECT 20.224 5.004 20.256 5.748 ;
  LAYER M1 ;
        RECT 20.224 5.844 20.256 6.084 ;
  LAYER M1 ;
        RECT 20.224 6.18 20.256 6.924 ;
  LAYER M1 ;
        RECT 20.224 7.02 20.256 7.26 ;
  LAYER M1 ;
        RECT 20.224 7.356 20.256 8.1 ;
  LAYER M1 ;
        RECT 20.224 8.196 20.256 8.436 ;
  LAYER M1 ;
        RECT 20.224 8.7 20.256 8.94 ;
  LAYER M1 ;
        RECT 20.304 0.3 20.336 1.044 ;
  LAYER M1 ;
        RECT 20.304 1.476 20.336 2.22 ;
  LAYER M1 ;
        RECT 20.304 2.652 20.336 3.396 ;
  LAYER M1 ;
        RECT 20.304 3.828 20.336 4.572 ;
  LAYER M1 ;
        RECT 20.304 5.004 20.336 5.748 ;
  LAYER M1 ;
        RECT 20.304 6.18 20.336 6.924 ;
  LAYER M1 ;
        RECT 20.304 7.356 20.336 8.1 ;
  LAYER M1 ;
        RECT 20.384 0.3 20.416 1.044 ;
  LAYER M1 ;
        RECT 20.384 1.14 20.416 1.38 ;
  LAYER M1 ;
        RECT 20.384 1.476 20.416 2.22 ;
  LAYER M1 ;
        RECT 20.384 2.316 20.416 2.556 ;
  LAYER M1 ;
        RECT 20.384 2.652 20.416 3.396 ;
  LAYER M1 ;
        RECT 20.384 3.492 20.416 3.732 ;
  LAYER M1 ;
        RECT 20.384 3.828 20.416 4.572 ;
  LAYER M1 ;
        RECT 20.384 4.668 20.416 4.908 ;
  LAYER M1 ;
        RECT 20.384 5.004 20.416 5.748 ;
  LAYER M1 ;
        RECT 20.384 5.844 20.416 6.084 ;
  LAYER M1 ;
        RECT 20.384 6.18 20.416 6.924 ;
  LAYER M1 ;
        RECT 20.384 7.02 20.416 7.26 ;
  LAYER M1 ;
        RECT 20.384 7.356 20.416 8.1 ;
  LAYER M1 ;
        RECT 20.384 8.196 20.416 8.436 ;
  LAYER M1 ;
        RECT 20.384 8.7 20.416 8.94 ;
  LAYER M1 ;
        RECT 20.464 0.3 20.496 1.044 ;
  LAYER M1 ;
        RECT 20.464 1.476 20.496 2.22 ;
  LAYER M1 ;
        RECT 20.464 2.652 20.496 3.396 ;
  LAYER M1 ;
        RECT 20.464 3.828 20.496 4.572 ;
  LAYER M1 ;
        RECT 20.464 5.004 20.496 5.748 ;
  LAYER M1 ;
        RECT 20.464 6.18 20.496 6.924 ;
  LAYER M1 ;
        RECT 20.464 7.356 20.496 8.1 ;
  LAYER M2 ;
        RECT 16.604 0.32 20.516 0.352 ;
  LAYER M2 ;
        RECT 16.684 0.404 20.436 0.436 ;
  LAYER M2 ;
        RECT 16.684 1.16 20.436 1.192 ;
  LAYER M2 ;
        RECT 16.844 0.488 20.276 0.52 ;
  LAYER M2 ;
        RECT 16.604 1.496 20.516 1.528 ;
  LAYER M2 ;
        RECT 16.844 1.58 20.276 1.612 ;
  LAYER M2 ;
        RECT 16.684 2.336 20.436 2.368 ;
  LAYER M2 ;
        RECT 16.684 1.664 20.436 1.696 ;
  LAYER M2 ;
        RECT 16.604 2.672 20.516 2.704 ;
  LAYER M2 ;
        RECT 16.684 2.756 20.436 2.788 ;
  LAYER M2 ;
        RECT 16.684 3.512 20.436 3.544 ;
  LAYER M2 ;
        RECT 16.844 2.84 20.276 2.872 ;
  LAYER M2 ;
        RECT 16.604 3.848 20.516 3.88 ;
  LAYER M2 ;
        RECT 16.844 3.932 20.276 3.964 ;
  LAYER M2 ;
        RECT 16.684 4.688 20.436 4.72 ;
  LAYER M2 ;
        RECT 16.684 4.016 20.436 4.048 ;
  LAYER M2 ;
        RECT 16.604 5.024 20.516 5.056 ;
  LAYER M2 ;
        RECT 16.684 5.108 20.436 5.14 ;
  LAYER M2 ;
        RECT 16.684 5.864 20.436 5.896 ;
  LAYER M2 ;
        RECT 16.844 5.192 20.276 5.224 ;
  LAYER M2 ;
        RECT 16.604 6.2 20.516 6.232 ;
  LAYER M2 ;
        RECT 16.844 6.284 20.276 6.316 ;
  LAYER M2 ;
        RECT 16.684 7.04 20.436 7.072 ;
  LAYER M2 ;
        RECT 16.684 6.368 20.436 6.4 ;
  LAYER M2 ;
        RECT 16.604 7.376 20.516 7.408 ;
  LAYER M2 ;
        RECT 16.684 7.46 20.436 7.492 ;
  LAYER M2 ;
        RECT 16.684 8.216 20.436 8.248 ;
  LAYER M2 ;
        RECT 16.844 7.544 20.276 7.576 ;
  LAYER M1 ;
        RECT 7.424 9.54 7.456 10.284 ;
  LAYER M1 ;
        RECT 7.424 10.38 7.456 10.62 ;
  LAYER M1 ;
        RECT 7.424 10.716 7.456 11.46 ;
  LAYER M1 ;
        RECT 7.424 11.556 7.456 11.796 ;
  LAYER M1 ;
        RECT 7.424 11.892 7.456 12.636 ;
  LAYER M1 ;
        RECT 7.424 12.732 7.456 12.972 ;
  LAYER M1 ;
        RECT 7.424 13.068 7.456 13.812 ;
  LAYER M1 ;
        RECT 7.424 13.908 7.456 14.148 ;
  LAYER M1 ;
        RECT 7.424 14.244 7.456 14.988 ;
  LAYER M1 ;
        RECT 7.424 15.084 7.456 15.324 ;
  LAYER M1 ;
        RECT 7.424 15.42 7.456 16.164 ;
  LAYER M1 ;
        RECT 7.424 16.26 7.456 16.5 ;
  LAYER M1 ;
        RECT 7.424 16.596 7.456 17.34 ;
  LAYER M1 ;
        RECT 7.424 17.436 7.456 17.676 ;
  LAYER M1 ;
        RECT 7.424 17.94 7.456 18.18 ;
  LAYER M1 ;
        RECT 7.344 9.54 7.376 10.284 ;
  LAYER M1 ;
        RECT 7.344 10.716 7.376 11.46 ;
  LAYER M1 ;
        RECT 7.344 11.892 7.376 12.636 ;
  LAYER M1 ;
        RECT 7.344 13.068 7.376 13.812 ;
  LAYER M1 ;
        RECT 7.344 14.244 7.376 14.988 ;
  LAYER M1 ;
        RECT 7.344 15.42 7.376 16.164 ;
  LAYER M1 ;
        RECT 7.344 16.596 7.376 17.34 ;
  LAYER M1 ;
        RECT 7.504 9.54 7.536 10.284 ;
  LAYER M1 ;
        RECT 7.504 10.716 7.536 11.46 ;
  LAYER M1 ;
        RECT 7.504 11.892 7.536 12.636 ;
  LAYER M1 ;
        RECT 7.504 13.068 7.536 13.812 ;
  LAYER M1 ;
        RECT 7.504 14.244 7.536 14.988 ;
  LAYER M1 ;
        RECT 7.504 15.42 7.536 16.164 ;
  LAYER M1 ;
        RECT 7.504 16.596 7.536 17.34 ;
  LAYER M1 ;
        RECT 7.584 9.54 7.616 10.284 ;
  LAYER M1 ;
        RECT 7.584 10.38 7.616 10.62 ;
  LAYER M1 ;
        RECT 7.584 10.716 7.616 11.46 ;
  LAYER M1 ;
        RECT 7.584 11.556 7.616 11.796 ;
  LAYER M1 ;
        RECT 7.584 11.892 7.616 12.636 ;
  LAYER M1 ;
        RECT 7.584 12.732 7.616 12.972 ;
  LAYER M1 ;
        RECT 7.584 13.068 7.616 13.812 ;
  LAYER M1 ;
        RECT 7.584 13.908 7.616 14.148 ;
  LAYER M1 ;
        RECT 7.584 14.244 7.616 14.988 ;
  LAYER M1 ;
        RECT 7.584 15.084 7.616 15.324 ;
  LAYER M1 ;
        RECT 7.584 15.42 7.616 16.164 ;
  LAYER M1 ;
        RECT 7.584 16.26 7.616 16.5 ;
  LAYER M1 ;
        RECT 7.584 16.596 7.616 17.34 ;
  LAYER M1 ;
        RECT 7.584 17.436 7.616 17.676 ;
  LAYER M1 ;
        RECT 7.584 17.94 7.616 18.18 ;
  LAYER M1 ;
        RECT 7.664 9.54 7.696 10.284 ;
  LAYER M1 ;
        RECT 7.664 10.716 7.696 11.46 ;
  LAYER M1 ;
        RECT 7.664 11.892 7.696 12.636 ;
  LAYER M1 ;
        RECT 7.664 13.068 7.696 13.812 ;
  LAYER M1 ;
        RECT 7.664 14.244 7.696 14.988 ;
  LAYER M1 ;
        RECT 7.664 15.42 7.696 16.164 ;
  LAYER M1 ;
        RECT 7.664 16.596 7.696 17.34 ;
  LAYER M1 ;
        RECT 7.744 9.54 7.776 10.284 ;
  LAYER M1 ;
        RECT 7.744 10.38 7.776 10.62 ;
  LAYER M1 ;
        RECT 7.744 10.716 7.776 11.46 ;
  LAYER M1 ;
        RECT 7.744 11.556 7.776 11.796 ;
  LAYER M1 ;
        RECT 7.744 11.892 7.776 12.636 ;
  LAYER M1 ;
        RECT 7.744 12.732 7.776 12.972 ;
  LAYER M1 ;
        RECT 7.744 13.068 7.776 13.812 ;
  LAYER M1 ;
        RECT 7.744 13.908 7.776 14.148 ;
  LAYER M1 ;
        RECT 7.744 14.244 7.776 14.988 ;
  LAYER M1 ;
        RECT 7.744 15.084 7.776 15.324 ;
  LAYER M1 ;
        RECT 7.744 15.42 7.776 16.164 ;
  LAYER M1 ;
        RECT 7.744 16.26 7.776 16.5 ;
  LAYER M1 ;
        RECT 7.744 16.596 7.776 17.34 ;
  LAYER M1 ;
        RECT 7.744 17.436 7.776 17.676 ;
  LAYER M1 ;
        RECT 7.744 17.94 7.776 18.18 ;
  LAYER M1 ;
        RECT 7.824 9.54 7.856 10.284 ;
  LAYER M1 ;
        RECT 7.824 10.716 7.856 11.46 ;
  LAYER M1 ;
        RECT 7.824 11.892 7.856 12.636 ;
  LAYER M1 ;
        RECT 7.824 13.068 7.856 13.812 ;
  LAYER M1 ;
        RECT 7.824 14.244 7.856 14.988 ;
  LAYER M1 ;
        RECT 7.824 15.42 7.856 16.164 ;
  LAYER M1 ;
        RECT 7.824 16.596 7.856 17.34 ;
  LAYER M1 ;
        RECT 7.904 9.54 7.936 10.284 ;
  LAYER M1 ;
        RECT 7.904 10.38 7.936 10.62 ;
  LAYER M1 ;
        RECT 7.904 10.716 7.936 11.46 ;
  LAYER M1 ;
        RECT 7.904 11.556 7.936 11.796 ;
  LAYER M1 ;
        RECT 7.904 11.892 7.936 12.636 ;
  LAYER M1 ;
        RECT 7.904 12.732 7.936 12.972 ;
  LAYER M1 ;
        RECT 7.904 13.068 7.936 13.812 ;
  LAYER M1 ;
        RECT 7.904 13.908 7.936 14.148 ;
  LAYER M1 ;
        RECT 7.904 14.244 7.936 14.988 ;
  LAYER M1 ;
        RECT 7.904 15.084 7.936 15.324 ;
  LAYER M1 ;
        RECT 7.904 15.42 7.936 16.164 ;
  LAYER M1 ;
        RECT 7.904 16.26 7.936 16.5 ;
  LAYER M1 ;
        RECT 7.904 16.596 7.936 17.34 ;
  LAYER M1 ;
        RECT 7.904 17.436 7.936 17.676 ;
  LAYER M1 ;
        RECT 7.904 17.94 7.936 18.18 ;
  LAYER M1 ;
        RECT 7.984 9.54 8.016 10.284 ;
  LAYER M1 ;
        RECT 7.984 10.716 8.016 11.46 ;
  LAYER M1 ;
        RECT 7.984 11.892 8.016 12.636 ;
  LAYER M1 ;
        RECT 7.984 13.068 8.016 13.812 ;
  LAYER M1 ;
        RECT 7.984 14.244 8.016 14.988 ;
  LAYER M1 ;
        RECT 7.984 15.42 8.016 16.164 ;
  LAYER M1 ;
        RECT 7.984 16.596 8.016 17.34 ;
  LAYER M1 ;
        RECT 8.064 9.54 8.096 10.284 ;
  LAYER M1 ;
        RECT 8.064 10.38 8.096 10.62 ;
  LAYER M1 ;
        RECT 8.064 10.716 8.096 11.46 ;
  LAYER M1 ;
        RECT 8.064 11.556 8.096 11.796 ;
  LAYER M1 ;
        RECT 8.064 11.892 8.096 12.636 ;
  LAYER M1 ;
        RECT 8.064 12.732 8.096 12.972 ;
  LAYER M1 ;
        RECT 8.064 13.068 8.096 13.812 ;
  LAYER M1 ;
        RECT 8.064 13.908 8.096 14.148 ;
  LAYER M1 ;
        RECT 8.064 14.244 8.096 14.988 ;
  LAYER M1 ;
        RECT 8.064 15.084 8.096 15.324 ;
  LAYER M1 ;
        RECT 8.064 15.42 8.096 16.164 ;
  LAYER M1 ;
        RECT 8.064 16.26 8.096 16.5 ;
  LAYER M1 ;
        RECT 8.064 16.596 8.096 17.34 ;
  LAYER M1 ;
        RECT 8.064 17.436 8.096 17.676 ;
  LAYER M1 ;
        RECT 8.064 17.94 8.096 18.18 ;
  LAYER M1 ;
        RECT 8.144 9.54 8.176 10.284 ;
  LAYER M1 ;
        RECT 8.144 10.716 8.176 11.46 ;
  LAYER M1 ;
        RECT 8.144 11.892 8.176 12.636 ;
  LAYER M1 ;
        RECT 8.144 13.068 8.176 13.812 ;
  LAYER M1 ;
        RECT 8.144 14.244 8.176 14.988 ;
  LAYER M1 ;
        RECT 8.144 15.42 8.176 16.164 ;
  LAYER M1 ;
        RECT 8.144 16.596 8.176 17.34 ;
  LAYER M1 ;
        RECT 8.224 9.54 8.256 10.284 ;
  LAYER M1 ;
        RECT 8.224 10.38 8.256 10.62 ;
  LAYER M1 ;
        RECT 8.224 10.716 8.256 11.46 ;
  LAYER M1 ;
        RECT 8.224 11.556 8.256 11.796 ;
  LAYER M1 ;
        RECT 8.224 11.892 8.256 12.636 ;
  LAYER M1 ;
        RECT 8.224 12.732 8.256 12.972 ;
  LAYER M1 ;
        RECT 8.224 13.068 8.256 13.812 ;
  LAYER M1 ;
        RECT 8.224 13.908 8.256 14.148 ;
  LAYER M1 ;
        RECT 8.224 14.244 8.256 14.988 ;
  LAYER M1 ;
        RECT 8.224 15.084 8.256 15.324 ;
  LAYER M1 ;
        RECT 8.224 15.42 8.256 16.164 ;
  LAYER M1 ;
        RECT 8.224 16.26 8.256 16.5 ;
  LAYER M1 ;
        RECT 8.224 16.596 8.256 17.34 ;
  LAYER M1 ;
        RECT 8.224 17.436 8.256 17.676 ;
  LAYER M1 ;
        RECT 8.224 17.94 8.256 18.18 ;
  LAYER M1 ;
        RECT 8.304 9.54 8.336 10.284 ;
  LAYER M1 ;
        RECT 8.304 10.716 8.336 11.46 ;
  LAYER M1 ;
        RECT 8.304 11.892 8.336 12.636 ;
  LAYER M1 ;
        RECT 8.304 13.068 8.336 13.812 ;
  LAYER M1 ;
        RECT 8.304 14.244 8.336 14.988 ;
  LAYER M1 ;
        RECT 8.304 15.42 8.336 16.164 ;
  LAYER M1 ;
        RECT 8.304 16.596 8.336 17.34 ;
  LAYER M1 ;
        RECT 8.384 9.54 8.416 10.284 ;
  LAYER M1 ;
        RECT 8.384 10.38 8.416 10.62 ;
  LAYER M1 ;
        RECT 8.384 10.716 8.416 11.46 ;
  LAYER M1 ;
        RECT 8.384 11.556 8.416 11.796 ;
  LAYER M1 ;
        RECT 8.384 11.892 8.416 12.636 ;
  LAYER M1 ;
        RECT 8.384 12.732 8.416 12.972 ;
  LAYER M1 ;
        RECT 8.384 13.068 8.416 13.812 ;
  LAYER M1 ;
        RECT 8.384 13.908 8.416 14.148 ;
  LAYER M1 ;
        RECT 8.384 14.244 8.416 14.988 ;
  LAYER M1 ;
        RECT 8.384 15.084 8.416 15.324 ;
  LAYER M1 ;
        RECT 8.384 15.42 8.416 16.164 ;
  LAYER M1 ;
        RECT 8.384 16.26 8.416 16.5 ;
  LAYER M1 ;
        RECT 8.384 16.596 8.416 17.34 ;
  LAYER M1 ;
        RECT 8.384 17.436 8.416 17.676 ;
  LAYER M1 ;
        RECT 8.384 17.94 8.416 18.18 ;
  LAYER M1 ;
        RECT 8.464 9.54 8.496 10.284 ;
  LAYER M1 ;
        RECT 8.464 10.716 8.496 11.46 ;
  LAYER M1 ;
        RECT 8.464 11.892 8.496 12.636 ;
  LAYER M1 ;
        RECT 8.464 13.068 8.496 13.812 ;
  LAYER M1 ;
        RECT 8.464 14.244 8.496 14.988 ;
  LAYER M1 ;
        RECT 8.464 15.42 8.496 16.164 ;
  LAYER M1 ;
        RECT 8.464 16.596 8.496 17.34 ;
  LAYER M1 ;
        RECT 8.544 9.54 8.576 10.284 ;
  LAYER M1 ;
        RECT 8.544 10.38 8.576 10.62 ;
  LAYER M1 ;
        RECT 8.544 10.716 8.576 11.46 ;
  LAYER M1 ;
        RECT 8.544 11.556 8.576 11.796 ;
  LAYER M1 ;
        RECT 8.544 11.892 8.576 12.636 ;
  LAYER M1 ;
        RECT 8.544 12.732 8.576 12.972 ;
  LAYER M1 ;
        RECT 8.544 13.068 8.576 13.812 ;
  LAYER M1 ;
        RECT 8.544 13.908 8.576 14.148 ;
  LAYER M1 ;
        RECT 8.544 14.244 8.576 14.988 ;
  LAYER M1 ;
        RECT 8.544 15.084 8.576 15.324 ;
  LAYER M1 ;
        RECT 8.544 15.42 8.576 16.164 ;
  LAYER M1 ;
        RECT 8.544 16.26 8.576 16.5 ;
  LAYER M1 ;
        RECT 8.544 16.596 8.576 17.34 ;
  LAYER M1 ;
        RECT 8.544 17.436 8.576 17.676 ;
  LAYER M1 ;
        RECT 8.544 17.94 8.576 18.18 ;
  LAYER M1 ;
        RECT 8.624 9.54 8.656 10.284 ;
  LAYER M1 ;
        RECT 8.624 10.716 8.656 11.46 ;
  LAYER M1 ;
        RECT 8.624 11.892 8.656 12.636 ;
  LAYER M1 ;
        RECT 8.624 13.068 8.656 13.812 ;
  LAYER M1 ;
        RECT 8.624 14.244 8.656 14.988 ;
  LAYER M1 ;
        RECT 8.624 15.42 8.656 16.164 ;
  LAYER M1 ;
        RECT 8.624 16.596 8.656 17.34 ;
  LAYER M1 ;
        RECT 8.704 9.54 8.736 10.284 ;
  LAYER M1 ;
        RECT 8.704 10.38 8.736 10.62 ;
  LAYER M1 ;
        RECT 8.704 10.716 8.736 11.46 ;
  LAYER M1 ;
        RECT 8.704 11.556 8.736 11.796 ;
  LAYER M1 ;
        RECT 8.704 11.892 8.736 12.636 ;
  LAYER M1 ;
        RECT 8.704 12.732 8.736 12.972 ;
  LAYER M1 ;
        RECT 8.704 13.068 8.736 13.812 ;
  LAYER M1 ;
        RECT 8.704 13.908 8.736 14.148 ;
  LAYER M1 ;
        RECT 8.704 14.244 8.736 14.988 ;
  LAYER M1 ;
        RECT 8.704 15.084 8.736 15.324 ;
  LAYER M1 ;
        RECT 8.704 15.42 8.736 16.164 ;
  LAYER M1 ;
        RECT 8.704 16.26 8.736 16.5 ;
  LAYER M1 ;
        RECT 8.704 16.596 8.736 17.34 ;
  LAYER M1 ;
        RECT 8.704 17.436 8.736 17.676 ;
  LAYER M1 ;
        RECT 8.704 17.94 8.736 18.18 ;
  LAYER M1 ;
        RECT 8.784 9.54 8.816 10.284 ;
  LAYER M1 ;
        RECT 8.784 10.716 8.816 11.46 ;
  LAYER M1 ;
        RECT 8.784 11.892 8.816 12.636 ;
  LAYER M1 ;
        RECT 8.784 13.068 8.816 13.812 ;
  LAYER M1 ;
        RECT 8.784 14.244 8.816 14.988 ;
  LAYER M1 ;
        RECT 8.784 15.42 8.816 16.164 ;
  LAYER M1 ;
        RECT 8.784 16.596 8.816 17.34 ;
  LAYER M1 ;
        RECT 8.864 9.54 8.896 10.284 ;
  LAYER M1 ;
        RECT 8.864 10.38 8.896 10.62 ;
  LAYER M1 ;
        RECT 8.864 10.716 8.896 11.46 ;
  LAYER M1 ;
        RECT 8.864 11.556 8.896 11.796 ;
  LAYER M1 ;
        RECT 8.864 11.892 8.896 12.636 ;
  LAYER M1 ;
        RECT 8.864 12.732 8.896 12.972 ;
  LAYER M1 ;
        RECT 8.864 13.068 8.896 13.812 ;
  LAYER M1 ;
        RECT 8.864 13.908 8.896 14.148 ;
  LAYER M1 ;
        RECT 8.864 14.244 8.896 14.988 ;
  LAYER M1 ;
        RECT 8.864 15.084 8.896 15.324 ;
  LAYER M1 ;
        RECT 8.864 15.42 8.896 16.164 ;
  LAYER M1 ;
        RECT 8.864 16.26 8.896 16.5 ;
  LAYER M1 ;
        RECT 8.864 16.596 8.896 17.34 ;
  LAYER M1 ;
        RECT 8.864 17.436 8.896 17.676 ;
  LAYER M1 ;
        RECT 8.864 17.94 8.896 18.18 ;
  LAYER M1 ;
        RECT 8.944 9.54 8.976 10.284 ;
  LAYER M1 ;
        RECT 8.944 10.716 8.976 11.46 ;
  LAYER M1 ;
        RECT 8.944 11.892 8.976 12.636 ;
  LAYER M1 ;
        RECT 8.944 13.068 8.976 13.812 ;
  LAYER M1 ;
        RECT 8.944 14.244 8.976 14.988 ;
  LAYER M1 ;
        RECT 8.944 15.42 8.976 16.164 ;
  LAYER M1 ;
        RECT 8.944 16.596 8.976 17.34 ;
  LAYER M1 ;
        RECT 9.024 9.54 9.056 10.284 ;
  LAYER M1 ;
        RECT 9.024 10.38 9.056 10.62 ;
  LAYER M1 ;
        RECT 9.024 10.716 9.056 11.46 ;
  LAYER M1 ;
        RECT 9.024 11.556 9.056 11.796 ;
  LAYER M1 ;
        RECT 9.024 11.892 9.056 12.636 ;
  LAYER M1 ;
        RECT 9.024 12.732 9.056 12.972 ;
  LAYER M1 ;
        RECT 9.024 13.068 9.056 13.812 ;
  LAYER M1 ;
        RECT 9.024 13.908 9.056 14.148 ;
  LAYER M1 ;
        RECT 9.024 14.244 9.056 14.988 ;
  LAYER M1 ;
        RECT 9.024 15.084 9.056 15.324 ;
  LAYER M1 ;
        RECT 9.024 15.42 9.056 16.164 ;
  LAYER M1 ;
        RECT 9.024 16.26 9.056 16.5 ;
  LAYER M1 ;
        RECT 9.024 16.596 9.056 17.34 ;
  LAYER M1 ;
        RECT 9.024 17.436 9.056 17.676 ;
  LAYER M1 ;
        RECT 9.024 17.94 9.056 18.18 ;
  LAYER M1 ;
        RECT 9.104 9.54 9.136 10.284 ;
  LAYER M1 ;
        RECT 9.104 10.716 9.136 11.46 ;
  LAYER M1 ;
        RECT 9.104 11.892 9.136 12.636 ;
  LAYER M1 ;
        RECT 9.104 13.068 9.136 13.812 ;
  LAYER M1 ;
        RECT 9.104 14.244 9.136 14.988 ;
  LAYER M1 ;
        RECT 9.104 15.42 9.136 16.164 ;
  LAYER M1 ;
        RECT 9.104 16.596 9.136 17.34 ;
  LAYER M1 ;
        RECT 9.184 9.54 9.216 10.284 ;
  LAYER M1 ;
        RECT 9.184 10.38 9.216 10.62 ;
  LAYER M1 ;
        RECT 9.184 10.716 9.216 11.46 ;
  LAYER M1 ;
        RECT 9.184 11.556 9.216 11.796 ;
  LAYER M1 ;
        RECT 9.184 11.892 9.216 12.636 ;
  LAYER M1 ;
        RECT 9.184 12.732 9.216 12.972 ;
  LAYER M1 ;
        RECT 9.184 13.068 9.216 13.812 ;
  LAYER M1 ;
        RECT 9.184 13.908 9.216 14.148 ;
  LAYER M1 ;
        RECT 9.184 14.244 9.216 14.988 ;
  LAYER M1 ;
        RECT 9.184 15.084 9.216 15.324 ;
  LAYER M1 ;
        RECT 9.184 15.42 9.216 16.164 ;
  LAYER M1 ;
        RECT 9.184 16.26 9.216 16.5 ;
  LAYER M1 ;
        RECT 9.184 16.596 9.216 17.34 ;
  LAYER M1 ;
        RECT 9.184 17.436 9.216 17.676 ;
  LAYER M1 ;
        RECT 9.184 17.94 9.216 18.18 ;
  LAYER M1 ;
        RECT 9.264 9.54 9.296 10.284 ;
  LAYER M1 ;
        RECT 9.264 10.716 9.296 11.46 ;
  LAYER M1 ;
        RECT 9.264 11.892 9.296 12.636 ;
  LAYER M1 ;
        RECT 9.264 13.068 9.296 13.812 ;
  LAYER M1 ;
        RECT 9.264 14.244 9.296 14.988 ;
  LAYER M1 ;
        RECT 9.264 15.42 9.296 16.164 ;
  LAYER M1 ;
        RECT 9.264 16.596 9.296 17.34 ;
  LAYER M2 ;
        RECT 7.324 9.56 9.316 9.592 ;
  LAYER M2 ;
        RECT 7.404 9.644 9.236 9.676 ;
  LAYER M2 ;
        RECT 7.404 10.4 9.236 10.432 ;
  LAYER M2 ;
        RECT 7.324 10.736 9.316 10.768 ;
  LAYER M2 ;
        RECT 7.404 10.82 9.236 10.852 ;
  LAYER M2 ;
        RECT 7.404 11.576 9.236 11.608 ;
  LAYER M2 ;
        RECT 7.324 11.912 9.316 11.944 ;
  LAYER M2 ;
        RECT 7.404 11.996 9.236 12.028 ;
  LAYER M2 ;
        RECT 7.404 12.752 9.236 12.784 ;
  LAYER M2 ;
        RECT 7.324 13.088 9.316 13.12 ;
  LAYER M2 ;
        RECT 7.404 13.172 9.236 13.204 ;
  LAYER M2 ;
        RECT 7.404 13.928 9.236 13.96 ;
  LAYER M2 ;
        RECT 7.324 14.264 9.316 14.296 ;
  LAYER M2 ;
        RECT 7.404 14.348 9.236 14.38 ;
  LAYER M2 ;
        RECT 7.404 15.104 9.236 15.136 ;
  LAYER M2 ;
        RECT 7.324 15.44 9.316 15.472 ;
  LAYER M2 ;
        RECT 7.404 15.524 9.236 15.556 ;
  LAYER M2 ;
        RECT 7.404 16.28 9.236 16.312 ;
  LAYER M2 ;
        RECT 7.324 16.616 9.316 16.648 ;
  LAYER M2 ;
        RECT 7.404 16.7 9.236 16.732 ;
  LAYER M2 ;
        RECT 7.404 17.456 9.236 17.488 ;
  LAYER M1 ;
        RECT 9.904 9.54 9.936 10.284 ;
  LAYER M1 ;
        RECT 9.904 10.38 9.936 10.62 ;
  LAYER M1 ;
        RECT 9.904 10.716 9.936 11.46 ;
  LAYER M1 ;
        RECT 9.904 11.556 9.936 11.796 ;
  LAYER M1 ;
        RECT 9.904 11.892 9.936 12.636 ;
  LAYER M1 ;
        RECT 9.904 12.732 9.936 12.972 ;
  LAYER M1 ;
        RECT 9.904 13.068 9.936 13.812 ;
  LAYER M1 ;
        RECT 9.904 13.908 9.936 14.148 ;
  LAYER M1 ;
        RECT 9.904 14.244 9.936 14.988 ;
  LAYER M1 ;
        RECT 9.904 15.084 9.936 15.324 ;
  LAYER M1 ;
        RECT 9.904 15.42 9.936 16.164 ;
  LAYER M1 ;
        RECT 9.904 16.26 9.936 16.5 ;
  LAYER M1 ;
        RECT 9.904 16.596 9.936 17.34 ;
  LAYER M1 ;
        RECT 9.904 17.436 9.936 17.676 ;
  LAYER M1 ;
        RECT 9.904 17.94 9.936 18.18 ;
  LAYER M1 ;
        RECT 9.824 9.54 9.856 10.284 ;
  LAYER M1 ;
        RECT 9.824 10.716 9.856 11.46 ;
  LAYER M1 ;
        RECT 9.824 11.892 9.856 12.636 ;
  LAYER M1 ;
        RECT 9.824 13.068 9.856 13.812 ;
  LAYER M1 ;
        RECT 9.824 14.244 9.856 14.988 ;
  LAYER M1 ;
        RECT 9.824 15.42 9.856 16.164 ;
  LAYER M1 ;
        RECT 9.824 16.596 9.856 17.34 ;
  LAYER M1 ;
        RECT 9.984 9.54 10.016 10.284 ;
  LAYER M1 ;
        RECT 9.984 10.716 10.016 11.46 ;
  LAYER M1 ;
        RECT 9.984 11.892 10.016 12.636 ;
  LAYER M1 ;
        RECT 9.984 13.068 10.016 13.812 ;
  LAYER M1 ;
        RECT 9.984 14.244 10.016 14.988 ;
  LAYER M1 ;
        RECT 9.984 15.42 10.016 16.164 ;
  LAYER M1 ;
        RECT 9.984 16.596 10.016 17.34 ;
  LAYER M1 ;
        RECT 10.544 9.54 10.576 10.284 ;
  LAYER M1 ;
        RECT 10.544 10.38 10.576 10.62 ;
  LAYER M1 ;
        RECT 10.544 10.716 10.576 11.46 ;
  LAYER M1 ;
        RECT 10.544 11.556 10.576 11.796 ;
  LAYER M1 ;
        RECT 10.544 11.892 10.576 12.636 ;
  LAYER M1 ;
        RECT 10.544 12.732 10.576 12.972 ;
  LAYER M1 ;
        RECT 10.544 13.068 10.576 13.812 ;
  LAYER M1 ;
        RECT 10.544 13.908 10.576 14.148 ;
  LAYER M1 ;
        RECT 10.544 14.244 10.576 14.988 ;
  LAYER M1 ;
        RECT 10.544 15.084 10.576 15.324 ;
  LAYER M1 ;
        RECT 10.544 15.42 10.576 16.164 ;
  LAYER M1 ;
        RECT 10.544 16.26 10.576 16.5 ;
  LAYER M1 ;
        RECT 10.544 16.596 10.576 17.34 ;
  LAYER M1 ;
        RECT 10.544 17.436 10.576 17.676 ;
  LAYER M1 ;
        RECT 10.544 17.94 10.576 18.18 ;
  LAYER M1 ;
        RECT 10.464 9.54 10.496 10.284 ;
  LAYER M1 ;
        RECT 10.464 10.716 10.496 11.46 ;
  LAYER M1 ;
        RECT 10.464 11.892 10.496 12.636 ;
  LAYER M1 ;
        RECT 10.464 13.068 10.496 13.812 ;
  LAYER M1 ;
        RECT 10.464 14.244 10.496 14.988 ;
  LAYER M1 ;
        RECT 10.464 15.42 10.496 16.164 ;
  LAYER M1 ;
        RECT 10.464 16.596 10.496 17.34 ;
  LAYER M1 ;
        RECT 10.624 9.54 10.656 10.284 ;
  LAYER M1 ;
        RECT 10.624 10.716 10.656 11.46 ;
  LAYER M1 ;
        RECT 10.624 11.892 10.656 12.636 ;
  LAYER M1 ;
        RECT 10.624 13.068 10.656 13.812 ;
  LAYER M1 ;
        RECT 10.624 14.244 10.656 14.988 ;
  LAYER M1 ;
        RECT 10.624 15.42 10.656 16.164 ;
  LAYER M1 ;
        RECT 10.624 16.596 10.656 17.34 ;
  LAYER M1 ;
        RECT 11.184 9.54 11.216 10.284 ;
  LAYER M1 ;
        RECT 11.184 10.38 11.216 10.62 ;
  LAYER M1 ;
        RECT 11.184 10.716 11.216 11.46 ;
  LAYER M1 ;
        RECT 11.184 11.556 11.216 11.796 ;
  LAYER M1 ;
        RECT 11.184 11.892 11.216 12.636 ;
  LAYER M1 ;
        RECT 11.184 12.732 11.216 12.972 ;
  LAYER M1 ;
        RECT 11.184 13.068 11.216 13.812 ;
  LAYER M1 ;
        RECT 11.184 13.908 11.216 14.148 ;
  LAYER M1 ;
        RECT 11.184 14.244 11.216 14.988 ;
  LAYER M1 ;
        RECT 11.184 15.084 11.216 15.324 ;
  LAYER M1 ;
        RECT 11.184 15.42 11.216 16.164 ;
  LAYER M1 ;
        RECT 11.184 16.26 11.216 16.5 ;
  LAYER M1 ;
        RECT 11.184 16.596 11.216 17.34 ;
  LAYER M1 ;
        RECT 11.184 17.436 11.216 17.676 ;
  LAYER M1 ;
        RECT 11.184 17.94 11.216 18.18 ;
  LAYER M1 ;
        RECT 11.104 9.54 11.136 10.284 ;
  LAYER M1 ;
        RECT 11.104 10.716 11.136 11.46 ;
  LAYER M1 ;
        RECT 11.104 11.892 11.136 12.636 ;
  LAYER M1 ;
        RECT 11.104 13.068 11.136 13.812 ;
  LAYER M1 ;
        RECT 11.104 14.244 11.136 14.988 ;
  LAYER M1 ;
        RECT 11.104 15.42 11.136 16.164 ;
  LAYER M1 ;
        RECT 11.104 16.596 11.136 17.34 ;
  LAYER M1 ;
        RECT 11.264 9.54 11.296 10.284 ;
  LAYER M1 ;
        RECT 11.264 10.716 11.296 11.46 ;
  LAYER M1 ;
        RECT 11.264 11.892 11.296 12.636 ;
  LAYER M1 ;
        RECT 11.264 13.068 11.296 13.812 ;
  LAYER M1 ;
        RECT 11.264 14.244 11.296 14.988 ;
  LAYER M1 ;
        RECT 11.264 15.42 11.296 16.164 ;
  LAYER M1 ;
        RECT 11.264 16.596 11.296 17.34 ;
  LAYER M1 ;
        RECT 11.824 9.54 11.856 10.284 ;
  LAYER M1 ;
        RECT 11.824 10.38 11.856 10.62 ;
  LAYER M1 ;
        RECT 11.824 10.716 11.856 11.46 ;
  LAYER M1 ;
        RECT 11.824 11.556 11.856 11.796 ;
  LAYER M1 ;
        RECT 11.824 11.892 11.856 12.636 ;
  LAYER M1 ;
        RECT 11.824 12.732 11.856 12.972 ;
  LAYER M1 ;
        RECT 11.824 13.068 11.856 13.812 ;
  LAYER M1 ;
        RECT 11.824 13.908 11.856 14.148 ;
  LAYER M1 ;
        RECT 11.824 14.244 11.856 14.988 ;
  LAYER M1 ;
        RECT 11.824 15.084 11.856 15.324 ;
  LAYER M1 ;
        RECT 11.824 15.42 11.856 16.164 ;
  LAYER M1 ;
        RECT 11.824 16.26 11.856 16.5 ;
  LAYER M1 ;
        RECT 11.824 16.596 11.856 17.34 ;
  LAYER M1 ;
        RECT 11.824 17.436 11.856 17.676 ;
  LAYER M1 ;
        RECT 11.824 17.94 11.856 18.18 ;
  LAYER M1 ;
        RECT 11.744 9.54 11.776 10.284 ;
  LAYER M1 ;
        RECT 11.744 10.716 11.776 11.46 ;
  LAYER M1 ;
        RECT 11.744 11.892 11.776 12.636 ;
  LAYER M1 ;
        RECT 11.744 13.068 11.776 13.812 ;
  LAYER M1 ;
        RECT 11.744 14.244 11.776 14.988 ;
  LAYER M1 ;
        RECT 11.744 15.42 11.776 16.164 ;
  LAYER M1 ;
        RECT 11.744 16.596 11.776 17.34 ;
  LAYER M1 ;
        RECT 11.904 9.54 11.936 10.284 ;
  LAYER M1 ;
        RECT 11.904 10.716 11.936 11.46 ;
  LAYER M1 ;
        RECT 11.904 11.892 11.936 12.636 ;
  LAYER M1 ;
        RECT 11.904 13.068 11.936 13.812 ;
  LAYER M1 ;
        RECT 11.904 14.244 11.936 14.988 ;
  LAYER M1 ;
        RECT 11.904 15.42 11.936 16.164 ;
  LAYER M1 ;
        RECT 11.904 16.596 11.936 17.34 ;
  LAYER M1 ;
        RECT 12.464 9.54 12.496 10.284 ;
  LAYER M1 ;
        RECT 12.464 10.38 12.496 10.62 ;
  LAYER M1 ;
        RECT 12.464 10.716 12.496 11.46 ;
  LAYER M1 ;
        RECT 12.464 11.556 12.496 11.796 ;
  LAYER M1 ;
        RECT 12.464 11.892 12.496 12.636 ;
  LAYER M1 ;
        RECT 12.464 12.732 12.496 12.972 ;
  LAYER M1 ;
        RECT 12.464 13.068 12.496 13.812 ;
  LAYER M1 ;
        RECT 12.464 13.908 12.496 14.148 ;
  LAYER M1 ;
        RECT 12.464 14.244 12.496 14.988 ;
  LAYER M1 ;
        RECT 12.464 15.084 12.496 15.324 ;
  LAYER M1 ;
        RECT 12.464 15.42 12.496 16.164 ;
  LAYER M1 ;
        RECT 12.464 16.26 12.496 16.5 ;
  LAYER M1 ;
        RECT 12.464 16.596 12.496 17.34 ;
  LAYER M1 ;
        RECT 12.464 17.436 12.496 17.676 ;
  LAYER M1 ;
        RECT 12.464 17.94 12.496 18.18 ;
  LAYER M1 ;
        RECT 12.384 9.54 12.416 10.284 ;
  LAYER M1 ;
        RECT 12.384 10.716 12.416 11.46 ;
  LAYER M1 ;
        RECT 12.384 11.892 12.416 12.636 ;
  LAYER M1 ;
        RECT 12.384 13.068 12.416 13.812 ;
  LAYER M1 ;
        RECT 12.384 14.244 12.416 14.988 ;
  LAYER M1 ;
        RECT 12.384 15.42 12.416 16.164 ;
  LAYER M1 ;
        RECT 12.384 16.596 12.416 17.34 ;
  LAYER M1 ;
        RECT 12.544 9.54 12.576 10.284 ;
  LAYER M1 ;
        RECT 12.544 10.716 12.576 11.46 ;
  LAYER M1 ;
        RECT 12.544 11.892 12.576 12.636 ;
  LAYER M1 ;
        RECT 12.544 13.068 12.576 13.812 ;
  LAYER M1 ;
        RECT 12.544 14.244 12.576 14.988 ;
  LAYER M1 ;
        RECT 12.544 15.42 12.576 16.164 ;
  LAYER M1 ;
        RECT 12.544 16.596 12.576 17.34 ;
  LAYER M1 ;
        RECT 13.104 9.54 13.136 10.284 ;
  LAYER M1 ;
        RECT 13.104 10.38 13.136 10.62 ;
  LAYER M1 ;
        RECT 13.104 10.716 13.136 11.46 ;
  LAYER M1 ;
        RECT 13.104 11.556 13.136 11.796 ;
  LAYER M1 ;
        RECT 13.104 11.892 13.136 12.636 ;
  LAYER M1 ;
        RECT 13.104 12.732 13.136 12.972 ;
  LAYER M1 ;
        RECT 13.104 13.068 13.136 13.812 ;
  LAYER M1 ;
        RECT 13.104 13.908 13.136 14.148 ;
  LAYER M1 ;
        RECT 13.104 14.244 13.136 14.988 ;
  LAYER M1 ;
        RECT 13.104 15.084 13.136 15.324 ;
  LAYER M1 ;
        RECT 13.104 15.42 13.136 16.164 ;
  LAYER M1 ;
        RECT 13.104 16.26 13.136 16.5 ;
  LAYER M1 ;
        RECT 13.104 16.596 13.136 17.34 ;
  LAYER M1 ;
        RECT 13.104 17.436 13.136 17.676 ;
  LAYER M1 ;
        RECT 13.104 17.94 13.136 18.18 ;
  LAYER M1 ;
        RECT 13.024 9.54 13.056 10.284 ;
  LAYER M1 ;
        RECT 13.024 10.716 13.056 11.46 ;
  LAYER M1 ;
        RECT 13.024 11.892 13.056 12.636 ;
  LAYER M1 ;
        RECT 13.024 13.068 13.056 13.812 ;
  LAYER M1 ;
        RECT 13.024 14.244 13.056 14.988 ;
  LAYER M1 ;
        RECT 13.024 15.42 13.056 16.164 ;
  LAYER M1 ;
        RECT 13.024 16.596 13.056 17.34 ;
  LAYER M1 ;
        RECT 13.184 9.54 13.216 10.284 ;
  LAYER M1 ;
        RECT 13.184 10.716 13.216 11.46 ;
  LAYER M1 ;
        RECT 13.184 11.892 13.216 12.636 ;
  LAYER M1 ;
        RECT 13.184 13.068 13.216 13.812 ;
  LAYER M1 ;
        RECT 13.184 14.244 13.216 14.988 ;
  LAYER M1 ;
        RECT 13.184 15.42 13.216 16.164 ;
  LAYER M1 ;
        RECT 13.184 16.596 13.216 17.34 ;
  LAYER M1 ;
        RECT 13.744 9.54 13.776 10.284 ;
  LAYER M1 ;
        RECT 13.744 10.38 13.776 10.62 ;
  LAYER M1 ;
        RECT 13.744 10.716 13.776 11.46 ;
  LAYER M1 ;
        RECT 13.744 11.556 13.776 11.796 ;
  LAYER M1 ;
        RECT 13.744 11.892 13.776 12.636 ;
  LAYER M1 ;
        RECT 13.744 12.732 13.776 12.972 ;
  LAYER M1 ;
        RECT 13.744 13.068 13.776 13.812 ;
  LAYER M1 ;
        RECT 13.744 13.908 13.776 14.148 ;
  LAYER M1 ;
        RECT 13.744 14.244 13.776 14.988 ;
  LAYER M1 ;
        RECT 13.744 15.084 13.776 15.324 ;
  LAYER M1 ;
        RECT 13.744 15.42 13.776 16.164 ;
  LAYER M1 ;
        RECT 13.744 16.26 13.776 16.5 ;
  LAYER M1 ;
        RECT 13.744 16.596 13.776 17.34 ;
  LAYER M1 ;
        RECT 13.744 17.436 13.776 17.676 ;
  LAYER M1 ;
        RECT 13.744 17.94 13.776 18.18 ;
  LAYER M1 ;
        RECT 13.664 9.54 13.696 10.284 ;
  LAYER M1 ;
        RECT 13.664 10.716 13.696 11.46 ;
  LAYER M1 ;
        RECT 13.664 11.892 13.696 12.636 ;
  LAYER M1 ;
        RECT 13.664 13.068 13.696 13.812 ;
  LAYER M1 ;
        RECT 13.664 14.244 13.696 14.988 ;
  LAYER M1 ;
        RECT 13.664 15.42 13.696 16.164 ;
  LAYER M1 ;
        RECT 13.664 16.596 13.696 17.34 ;
  LAYER M1 ;
        RECT 13.824 9.54 13.856 10.284 ;
  LAYER M1 ;
        RECT 13.824 10.716 13.856 11.46 ;
  LAYER M1 ;
        RECT 13.824 11.892 13.856 12.636 ;
  LAYER M1 ;
        RECT 13.824 13.068 13.856 13.812 ;
  LAYER M1 ;
        RECT 13.824 14.244 13.856 14.988 ;
  LAYER M1 ;
        RECT 13.824 15.42 13.856 16.164 ;
  LAYER M1 ;
        RECT 13.824 16.596 13.856 17.34 ;
  LAYER M1 ;
        RECT 14.384 9.54 14.416 10.284 ;
  LAYER M1 ;
        RECT 14.384 10.38 14.416 10.62 ;
  LAYER M1 ;
        RECT 14.384 10.716 14.416 11.46 ;
  LAYER M1 ;
        RECT 14.384 11.556 14.416 11.796 ;
  LAYER M1 ;
        RECT 14.384 11.892 14.416 12.636 ;
  LAYER M1 ;
        RECT 14.384 12.732 14.416 12.972 ;
  LAYER M1 ;
        RECT 14.384 13.068 14.416 13.812 ;
  LAYER M1 ;
        RECT 14.384 13.908 14.416 14.148 ;
  LAYER M1 ;
        RECT 14.384 14.244 14.416 14.988 ;
  LAYER M1 ;
        RECT 14.384 15.084 14.416 15.324 ;
  LAYER M1 ;
        RECT 14.384 15.42 14.416 16.164 ;
  LAYER M1 ;
        RECT 14.384 16.26 14.416 16.5 ;
  LAYER M1 ;
        RECT 14.384 16.596 14.416 17.34 ;
  LAYER M1 ;
        RECT 14.384 17.436 14.416 17.676 ;
  LAYER M1 ;
        RECT 14.384 17.94 14.416 18.18 ;
  LAYER M1 ;
        RECT 14.304 9.54 14.336 10.284 ;
  LAYER M1 ;
        RECT 14.304 10.716 14.336 11.46 ;
  LAYER M1 ;
        RECT 14.304 11.892 14.336 12.636 ;
  LAYER M1 ;
        RECT 14.304 13.068 14.336 13.812 ;
  LAYER M1 ;
        RECT 14.304 14.244 14.336 14.988 ;
  LAYER M1 ;
        RECT 14.304 15.42 14.336 16.164 ;
  LAYER M1 ;
        RECT 14.304 16.596 14.336 17.34 ;
  LAYER M1 ;
        RECT 14.464 9.54 14.496 10.284 ;
  LAYER M1 ;
        RECT 14.464 10.716 14.496 11.46 ;
  LAYER M1 ;
        RECT 14.464 11.892 14.496 12.636 ;
  LAYER M1 ;
        RECT 14.464 13.068 14.496 13.812 ;
  LAYER M1 ;
        RECT 14.464 14.244 14.496 14.988 ;
  LAYER M1 ;
        RECT 14.464 15.42 14.496 16.164 ;
  LAYER M1 ;
        RECT 14.464 16.596 14.496 17.34 ;
  LAYER M1 ;
        RECT 15.024 9.54 15.056 10.284 ;
  LAYER M1 ;
        RECT 15.024 10.38 15.056 10.62 ;
  LAYER M1 ;
        RECT 15.024 10.716 15.056 11.46 ;
  LAYER M1 ;
        RECT 15.024 11.556 15.056 11.796 ;
  LAYER M1 ;
        RECT 15.024 11.892 15.056 12.636 ;
  LAYER M1 ;
        RECT 15.024 12.732 15.056 12.972 ;
  LAYER M1 ;
        RECT 15.024 13.068 15.056 13.812 ;
  LAYER M1 ;
        RECT 15.024 13.908 15.056 14.148 ;
  LAYER M1 ;
        RECT 15.024 14.244 15.056 14.988 ;
  LAYER M1 ;
        RECT 15.024 15.084 15.056 15.324 ;
  LAYER M1 ;
        RECT 15.024 15.42 15.056 16.164 ;
  LAYER M1 ;
        RECT 15.024 16.26 15.056 16.5 ;
  LAYER M1 ;
        RECT 15.024 16.596 15.056 17.34 ;
  LAYER M1 ;
        RECT 15.024 17.436 15.056 17.676 ;
  LAYER M1 ;
        RECT 15.024 17.94 15.056 18.18 ;
  LAYER M1 ;
        RECT 14.944 9.54 14.976 10.284 ;
  LAYER M1 ;
        RECT 14.944 10.716 14.976 11.46 ;
  LAYER M1 ;
        RECT 14.944 11.892 14.976 12.636 ;
  LAYER M1 ;
        RECT 14.944 13.068 14.976 13.812 ;
  LAYER M1 ;
        RECT 14.944 14.244 14.976 14.988 ;
  LAYER M1 ;
        RECT 14.944 15.42 14.976 16.164 ;
  LAYER M1 ;
        RECT 14.944 16.596 14.976 17.34 ;
  LAYER M1 ;
        RECT 15.104 9.54 15.136 10.284 ;
  LAYER M1 ;
        RECT 15.104 10.716 15.136 11.46 ;
  LAYER M1 ;
        RECT 15.104 11.892 15.136 12.636 ;
  LAYER M1 ;
        RECT 15.104 13.068 15.136 13.812 ;
  LAYER M1 ;
        RECT 15.104 14.244 15.136 14.988 ;
  LAYER M1 ;
        RECT 15.104 15.42 15.136 16.164 ;
  LAYER M1 ;
        RECT 15.104 16.596 15.136 17.34 ;
  LAYER M1 ;
        RECT 15.664 9.54 15.696 10.284 ;
  LAYER M1 ;
        RECT 15.664 10.38 15.696 10.62 ;
  LAYER M1 ;
        RECT 15.664 10.716 15.696 11.46 ;
  LAYER M1 ;
        RECT 15.664 11.556 15.696 11.796 ;
  LAYER M1 ;
        RECT 15.664 11.892 15.696 12.636 ;
  LAYER M1 ;
        RECT 15.664 12.732 15.696 12.972 ;
  LAYER M1 ;
        RECT 15.664 13.068 15.696 13.812 ;
  LAYER M1 ;
        RECT 15.664 13.908 15.696 14.148 ;
  LAYER M1 ;
        RECT 15.664 14.244 15.696 14.988 ;
  LAYER M1 ;
        RECT 15.664 15.084 15.696 15.324 ;
  LAYER M1 ;
        RECT 15.664 15.42 15.696 16.164 ;
  LAYER M1 ;
        RECT 15.664 16.26 15.696 16.5 ;
  LAYER M1 ;
        RECT 15.664 16.596 15.696 17.34 ;
  LAYER M1 ;
        RECT 15.664 17.436 15.696 17.676 ;
  LAYER M1 ;
        RECT 15.664 17.94 15.696 18.18 ;
  LAYER M1 ;
        RECT 15.584 9.54 15.616 10.284 ;
  LAYER M1 ;
        RECT 15.584 10.716 15.616 11.46 ;
  LAYER M1 ;
        RECT 15.584 11.892 15.616 12.636 ;
  LAYER M1 ;
        RECT 15.584 13.068 15.616 13.812 ;
  LAYER M1 ;
        RECT 15.584 14.244 15.616 14.988 ;
  LAYER M1 ;
        RECT 15.584 15.42 15.616 16.164 ;
  LAYER M1 ;
        RECT 15.584 16.596 15.616 17.34 ;
  LAYER M1 ;
        RECT 15.744 9.54 15.776 10.284 ;
  LAYER M1 ;
        RECT 15.744 10.716 15.776 11.46 ;
  LAYER M1 ;
        RECT 15.744 11.892 15.776 12.636 ;
  LAYER M1 ;
        RECT 15.744 13.068 15.776 13.812 ;
  LAYER M1 ;
        RECT 15.744 14.244 15.776 14.988 ;
  LAYER M1 ;
        RECT 15.744 15.42 15.776 16.164 ;
  LAYER M1 ;
        RECT 15.744 16.596 15.776 17.34 ;
  LAYER M1 ;
        RECT 16.304 9.54 16.336 10.284 ;
  LAYER M1 ;
        RECT 16.304 10.38 16.336 10.62 ;
  LAYER M1 ;
        RECT 16.304 10.716 16.336 11.46 ;
  LAYER M1 ;
        RECT 16.304 11.556 16.336 11.796 ;
  LAYER M1 ;
        RECT 16.304 11.892 16.336 12.636 ;
  LAYER M1 ;
        RECT 16.304 12.732 16.336 12.972 ;
  LAYER M1 ;
        RECT 16.304 13.068 16.336 13.812 ;
  LAYER M1 ;
        RECT 16.304 13.908 16.336 14.148 ;
  LAYER M1 ;
        RECT 16.304 14.244 16.336 14.988 ;
  LAYER M1 ;
        RECT 16.304 15.084 16.336 15.324 ;
  LAYER M1 ;
        RECT 16.304 15.42 16.336 16.164 ;
  LAYER M1 ;
        RECT 16.304 16.26 16.336 16.5 ;
  LAYER M1 ;
        RECT 16.304 16.596 16.336 17.34 ;
  LAYER M1 ;
        RECT 16.304 17.436 16.336 17.676 ;
  LAYER M1 ;
        RECT 16.304 17.94 16.336 18.18 ;
  LAYER M1 ;
        RECT 16.224 9.54 16.256 10.284 ;
  LAYER M1 ;
        RECT 16.224 10.716 16.256 11.46 ;
  LAYER M1 ;
        RECT 16.224 11.892 16.256 12.636 ;
  LAYER M1 ;
        RECT 16.224 13.068 16.256 13.812 ;
  LAYER M1 ;
        RECT 16.224 14.244 16.256 14.988 ;
  LAYER M1 ;
        RECT 16.224 15.42 16.256 16.164 ;
  LAYER M1 ;
        RECT 16.224 16.596 16.256 17.34 ;
  LAYER M1 ;
        RECT 16.384 9.54 16.416 10.284 ;
  LAYER M1 ;
        RECT 16.384 10.716 16.416 11.46 ;
  LAYER M1 ;
        RECT 16.384 11.892 16.416 12.636 ;
  LAYER M1 ;
        RECT 16.384 13.068 16.416 13.812 ;
  LAYER M1 ;
        RECT 16.384 14.244 16.416 14.988 ;
  LAYER M1 ;
        RECT 16.384 15.42 16.416 16.164 ;
  LAYER M1 ;
        RECT 16.384 16.596 16.416 17.34 ;
  LAYER M1 ;
        RECT 16.944 9.54 16.976 10.284 ;
  LAYER M1 ;
        RECT 16.944 10.38 16.976 10.62 ;
  LAYER M1 ;
        RECT 16.944 10.716 16.976 11.46 ;
  LAYER M1 ;
        RECT 16.944 11.556 16.976 11.796 ;
  LAYER M1 ;
        RECT 16.944 11.892 16.976 12.636 ;
  LAYER M1 ;
        RECT 16.944 12.732 16.976 12.972 ;
  LAYER M1 ;
        RECT 16.944 13.068 16.976 13.812 ;
  LAYER M1 ;
        RECT 16.944 13.908 16.976 14.148 ;
  LAYER M1 ;
        RECT 16.944 14.244 16.976 14.988 ;
  LAYER M1 ;
        RECT 16.944 15.084 16.976 15.324 ;
  LAYER M1 ;
        RECT 16.944 15.42 16.976 16.164 ;
  LAYER M1 ;
        RECT 16.944 16.26 16.976 16.5 ;
  LAYER M1 ;
        RECT 16.944 16.596 16.976 17.34 ;
  LAYER M1 ;
        RECT 16.944 17.436 16.976 17.676 ;
  LAYER M1 ;
        RECT 16.944 17.94 16.976 18.18 ;
  LAYER M1 ;
        RECT 16.864 9.54 16.896 10.284 ;
  LAYER M1 ;
        RECT 16.864 10.716 16.896 11.46 ;
  LAYER M1 ;
        RECT 16.864 11.892 16.896 12.636 ;
  LAYER M1 ;
        RECT 16.864 13.068 16.896 13.812 ;
  LAYER M1 ;
        RECT 16.864 14.244 16.896 14.988 ;
  LAYER M1 ;
        RECT 16.864 15.42 16.896 16.164 ;
  LAYER M1 ;
        RECT 16.864 16.596 16.896 17.34 ;
  LAYER M1 ;
        RECT 17.024 9.54 17.056 10.284 ;
  LAYER M1 ;
        RECT 17.024 10.716 17.056 11.46 ;
  LAYER M1 ;
        RECT 17.024 11.892 17.056 12.636 ;
  LAYER M1 ;
        RECT 17.024 13.068 17.056 13.812 ;
  LAYER M1 ;
        RECT 17.024 14.244 17.056 14.988 ;
  LAYER M1 ;
        RECT 17.024 15.42 17.056 16.164 ;
  LAYER M1 ;
        RECT 17.024 16.596 17.056 17.34 ;
  LAYER M1 ;
        RECT 17.584 9.54 17.616 10.284 ;
  LAYER M1 ;
        RECT 17.584 10.38 17.616 10.62 ;
  LAYER M1 ;
        RECT 17.584 10.716 17.616 11.46 ;
  LAYER M1 ;
        RECT 17.584 11.556 17.616 11.796 ;
  LAYER M1 ;
        RECT 17.584 11.892 17.616 12.636 ;
  LAYER M1 ;
        RECT 17.584 12.732 17.616 12.972 ;
  LAYER M1 ;
        RECT 17.584 13.068 17.616 13.812 ;
  LAYER M1 ;
        RECT 17.584 13.908 17.616 14.148 ;
  LAYER M1 ;
        RECT 17.584 14.244 17.616 14.988 ;
  LAYER M1 ;
        RECT 17.584 15.084 17.616 15.324 ;
  LAYER M1 ;
        RECT 17.584 15.42 17.616 16.164 ;
  LAYER M1 ;
        RECT 17.584 16.26 17.616 16.5 ;
  LAYER M1 ;
        RECT 17.584 16.596 17.616 17.34 ;
  LAYER M1 ;
        RECT 17.584 17.436 17.616 17.676 ;
  LAYER M1 ;
        RECT 17.584 17.94 17.616 18.18 ;
  LAYER M1 ;
        RECT 17.504 9.54 17.536 10.284 ;
  LAYER M1 ;
        RECT 17.504 10.716 17.536 11.46 ;
  LAYER M1 ;
        RECT 17.504 11.892 17.536 12.636 ;
  LAYER M1 ;
        RECT 17.504 13.068 17.536 13.812 ;
  LAYER M1 ;
        RECT 17.504 14.244 17.536 14.988 ;
  LAYER M1 ;
        RECT 17.504 15.42 17.536 16.164 ;
  LAYER M1 ;
        RECT 17.504 16.596 17.536 17.34 ;
  LAYER M1 ;
        RECT 17.664 9.54 17.696 10.284 ;
  LAYER M1 ;
        RECT 17.664 10.716 17.696 11.46 ;
  LAYER M1 ;
        RECT 17.664 11.892 17.696 12.636 ;
  LAYER M1 ;
        RECT 17.664 13.068 17.696 13.812 ;
  LAYER M1 ;
        RECT 17.664 14.244 17.696 14.988 ;
  LAYER M1 ;
        RECT 17.664 15.42 17.696 16.164 ;
  LAYER M1 ;
        RECT 17.664 16.596 17.696 17.34 ;
  LAYER M1 ;
        RECT 18.224 9.54 18.256 10.284 ;
  LAYER M1 ;
        RECT 18.224 10.38 18.256 10.62 ;
  LAYER M1 ;
        RECT 18.224 10.716 18.256 11.46 ;
  LAYER M1 ;
        RECT 18.224 11.556 18.256 11.796 ;
  LAYER M1 ;
        RECT 18.224 11.892 18.256 12.636 ;
  LAYER M1 ;
        RECT 18.224 12.732 18.256 12.972 ;
  LAYER M1 ;
        RECT 18.224 13.068 18.256 13.812 ;
  LAYER M1 ;
        RECT 18.224 13.908 18.256 14.148 ;
  LAYER M1 ;
        RECT 18.224 14.244 18.256 14.988 ;
  LAYER M1 ;
        RECT 18.224 15.084 18.256 15.324 ;
  LAYER M1 ;
        RECT 18.224 15.42 18.256 16.164 ;
  LAYER M1 ;
        RECT 18.224 16.26 18.256 16.5 ;
  LAYER M1 ;
        RECT 18.224 16.596 18.256 17.34 ;
  LAYER M1 ;
        RECT 18.224 17.436 18.256 17.676 ;
  LAYER M1 ;
        RECT 18.224 17.94 18.256 18.18 ;
  LAYER M1 ;
        RECT 18.144 9.54 18.176 10.284 ;
  LAYER M1 ;
        RECT 18.144 10.716 18.176 11.46 ;
  LAYER M1 ;
        RECT 18.144 11.892 18.176 12.636 ;
  LAYER M1 ;
        RECT 18.144 13.068 18.176 13.812 ;
  LAYER M1 ;
        RECT 18.144 14.244 18.176 14.988 ;
  LAYER M1 ;
        RECT 18.144 15.42 18.176 16.164 ;
  LAYER M1 ;
        RECT 18.144 16.596 18.176 17.34 ;
  LAYER M1 ;
        RECT 18.304 9.54 18.336 10.284 ;
  LAYER M1 ;
        RECT 18.304 10.716 18.336 11.46 ;
  LAYER M1 ;
        RECT 18.304 11.892 18.336 12.636 ;
  LAYER M1 ;
        RECT 18.304 13.068 18.336 13.812 ;
  LAYER M1 ;
        RECT 18.304 14.244 18.336 14.988 ;
  LAYER M1 ;
        RECT 18.304 15.42 18.336 16.164 ;
  LAYER M1 ;
        RECT 18.304 16.596 18.336 17.34 ;
  LAYER M1 ;
        RECT 18.864 9.54 18.896 10.284 ;
  LAYER M1 ;
        RECT 18.864 10.38 18.896 10.62 ;
  LAYER M1 ;
        RECT 18.864 10.716 18.896 11.46 ;
  LAYER M1 ;
        RECT 18.864 11.556 18.896 11.796 ;
  LAYER M1 ;
        RECT 18.864 11.892 18.896 12.636 ;
  LAYER M1 ;
        RECT 18.864 12.732 18.896 12.972 ;
  LAYER M1 ;
        RECT 18.864 13.068 18.896 13.812 ;
  LAYER M1 ;
        RECT 18.864 13.908 18.896 14.148 ;
  LAYER M1 ;
        RECT 18.864 14.244 18.896 14.988 ;
  LAYER M1 ;
        RECT 18.864 15.084 18.896 15.324 ;
  LAYER M1 ;
        RECT 18.864 15.42 18.896 16.164 ;
  LAYER M1 ;
        RECT 18.864 16.26 18.896 16.5 ;
  LAYER M1 ;
        RECT 18.864 16.596 18.896 17.34 ;
  LAYER M1 ;
        RECT 18.864 17.436 18.896 17.676 ;
  LAYER M1 ;
        RECT 18.864 17.94 18.896 18.18 ;
  LAYER M1 ;
        RECT 18.784 9.54 18.816 10.284 ;
  LAYER M1 ;
        RECT 18.784 10.716 18.816 11.46 ;
  LAYER M1 ;
        RECT 18.784 11.892 18.816 12.636 ;
  LAYER M1 ;
        RECT 18.784 13.068 18.816 13.812 ;
  LAYER M1 ;
        RECT 18.784 14.244 18.816 14.988 ;
  LAYER M1 ;
        RECT 18.784 15.42 18.816 16.164 ;
  LAYER M1 ;
        RECT 18.784 16.596 18.816 17.34 ;
  LAYER M1 ;
        RECT 18.944 9.54 18.976 10.284 ;
  LAYER M1 ;
        RECT 18.944 10.716 18.976 11.46 ;
  LAYER M1 ;
        RECT 18.944 11.892 18.976 12.636 ;
  LAYER M1 ;
        RECT 18.944 13.068 18.976 13.812 ;
  LAYER M1 ;
        RECT 18.944 14.244 18.976 14.988 ;
  LAYER M1 ;
        RECT 18.944 15.42 18.976 16.164 ;
  LAYER M1 ;
        RECT 18.944 16.596 18.976 17.34 ;
  LAYER M1 ;
        RECT 19.504 9.54 19.536 10.284 ;
  LAYER M1 ;
        RECT 19.504 10.38 19.536 10.62 ;
  LAYER M1 ;
        RECT 19.504 10.716 19.536 11.46 ;
  LAYER M1 ;
        RECT 19.504 11.556 19.536 11.796 ;
  LAYER M1 ;
        RECT 19.504 11.892 19.536 12.636 ;
  LAYER M1 ;
        RECT 19.504 12.732 19.536 12.972 ;
  LAYER M1 ;
        RECT 19.504 13.068 19.536 13.812 ;
  LAYER M1 ;
        RECT 19.504 13.908 19.536 14.148 ;
  LAYER M1 ;
        RECT 19.504 14.244 19.536 14.988 ;
  LAYER M1 ;
        RECT 19.504 15.084 19.536 15.324 ;
  LAYER M1 ;
        RECT 19.504 15.42 19.536 16.164 ;
  LAYER M1 ;
        RECT 19.504 16.26 19.536 16.5 ;
  LAYER M1 ;
        RECT 19.504 16.596 19.536 17.34 ;
  LAYER M1 ;
        RECT 19.504 17.436 19.536 17.676 ;
  LAYER M1 ;
        RECT 19.504 17.94 19.536 18.18 ;
  LAYER M1 ;
        RECT 19.424 9.54 19.456 10.284 ;
  LAYER M1 ;
        RECT 19.424 10.716 19.456 11.46 ;
  LAYER M1 ;
        RECT 19.424 11.892 19.456 12.636 ;
  LAYER M1 ;
        RECT 19.424 13.068 19.456 13.812 ;
  LAYER M1 ;
        RECT 19.424 14.244 19.456 14.988 ;
  LAYER M1 ;
        RECT 19.424 15.42 19.456 16.164 ;
  LAYER M1 ;
        RECT 19.424 16.596 19.456 17.34 ;
  LAYER M1 ;
        RECT 19.584 9.54 19.616 10.284 ;
  LAYER M1 ;
        RECT 19.584 10.716 19.616 11.46 ;
  LAYER M1 ;
        RECT 19.584 11.892 19.616 12.636 ;
  LAYER M1 ;
        RECT 19.584 13.068 19.616 13.812 ;
  LAYER M1 ;
        RECT 19.584 14.244 19.616 14.988 ;
  LAYER M1 ;
        RECT 19.584 15.42 19.616 16.164 ;
  LAYER M1 ;
        RECT 19.584 16.596 19.616 17.34 ;
  LAYER M1 ;
        RECT 20.144 9.54 20.176 10.284 ;
  LAYER M1 ;
        RECT 20.144 10.38 20.176 10.62 ;
  LAYER M1 ;
        RECT 20.144 10.716 20.176 11.46 ;
  LAYER M1 ;
        RECT 20.144 11.556 20.176 11.796 ;
  LAYER M1 ;
        RECT 20.144 11.892 20.176 12.636 ;
  LAYER M1 ;
        RECT 20.144 12.732 20.176 12.972 ;
  LAYER M1 ;
        RECT 20.144 13.068 20.176 13.812 ;
  LAYER M1 ;
        RECT 20.144 13.908 20.176 14.148 ;
  LAYER M1 ;
        RECT 20.144 14.244 20.176 14.988 ;
  LAYER M1 ;
        RECT 20.144 15.084 20.176 15.324 ;
  LAYER M1 ;
        RECT 20.144 15.42 20.176 16.164 ;
  LAYER M1 ;
        RECT 20.144 16.26 20.176 16.5 ;
  LAYER M1 ;
        RECT 20.144 16.596 20.176 17.34 ;
  LAYER M1 ;
        RECT 20.144 17.436 20.176 17.676 ;
  LAYER M1 ;
        RECT 20.144 17.94 20.176 18.18 ;
  LAYER M1 ;
        RECT 20.064 9.54 20.096 10.284 ;
  LAYER M1 ;
        RECT 20.064 10.716 20.096 11.46 ;
  LAYER M1 ;
        RECT 20.064 11.892 20.096 12.636 ;
  LAYER M1 ;
        RECT 20.064 13.068 20.096 13.812 ;
  LAYER M1 ;
        RECT 20.064 14.244 20.096 14.988 ;
  LAYER M1 ;
        RECT 20.064 15.42 20.096 16.164 ;
  LAYER M1 ;
        RECT 20.064 16.596 20.096 17.34 ;
  LAYER M1 ;
        RECT 20.224 9.54 20.256 10.284 ;
  LAYER M1 ;
        RECT 20.224 10.716 20.256 11.46 ;
  LAYER M1 ;
        RECT 20.224 11.892 20.256 12.636 ;
  LAYER M1 ;
        RECT 20.224 13.068 20.256 13.812 ;
  LAYER M1 ;
        RECT 20.224 14.244 20.256 14.988 ;
  LAYER M1 ;
        RECT 20.224 15.42 20.256 16.164 ;
  LAYER M1 ;
        RECT 20.224 16.596 20.256 17.34 ;
  LAYER M1 ;
        RECT 20.784 9.54 20.816 10.284 ;
  LAYER M1 ;
        RECT 20.784 10.38 20.816 10.62 ;
  LAYER M1 ;
        RECT 20.784 10.716 20.816 11.46 ;
  LAYER M1 ;
        RECT 20.784 11.556 20.816 11.796 ;
  LAYER M1 ;
        RECT 20.784 11.892 20.816 12.636 ;
  LAYER M1 ;
        RECT 20.784 12.732 20.816 12.972 ;
  LAYER M1 ;
        RECT 20.784 13.068 20.816 13.812 ;
  LAYER M1 ;
        RECT 20.784 13.908 20.816 14.148 ;
  LAYER M1 ;
        RECT 20.784 14.244 20.816 14.988 ;
  LAYER M1 ;
        RECT 20.784 15.084 20.816 15.324 ;
  LAYER M1 ;
        RECT 20.784 15.42 20.816 16.164 ;
  LAYER M1 ;
        RECT 20.784 16.26 20.816 16.5 ;
  LAYER M1 ;
        RECT 20.784 16.596 20.816 17.34 ;
  LAYER M1 ;
        RECT 20.784 17.436 20.816 17.676 ;
  LAYER M1 ;
        RECT 20.784 17.94 20.816 18.18 ;
  LAYER M1 ;
        RECT 20.704 9.54 20.736 10.284 ;
  LAYER M1 ;
        RECT 20.704 10.716 20.736 11.46 ;
  LAYER M1 ;
        RECT 20.704 11.892 20.736 12.636 ;
  LAYER M1 ;
        RECT 20.704 13.068 20.736 13.812 ;
  LAYER M1 ;
        RECT 20.704 14.244 20.736 14.988 ;
  LAYER M1 ;
        RECT 20.704 15.42 20.736 16.164 ;
  LAYER M1 ;
        RECT 20.704 16.596 20.736 17.34 ;
  LAYER M1 ;
        RECT 20.864 9.54 20.896 10.284 ;
  LAYER M1 ;
        RECT 20.864 10.716 20.896 11.46 ;
  LAYER M1 ;
        RECT 20.864 11.892 20.896 12.636 ;
  LAYER M1 ;
        RECT 20.864 13.068 20.896 13.812 ;
  LAYER M1 ;
        RECT 20.864 14.244 20.896 14.988 ;
  LAYER M1 ;
        RECT 20.864 15.42 20.896 16.164 ;
  LAYER M1 ;
        RECT 20.864 16.596 20.896 17.34 ;
  LAYER M1 ;
        RECT 21.424 9.54 21.456 10.284 ;
  LAYER M1 ;
        RECT 21.424 10.38 21.456 10.62 ;
  LAYER M1 ;
        RECT 21.424 10.716 21.456 11.46 ;
  LAYER M1 ;
        RECT 21.424 11.556 21.456 11.796 ;
  LAYER M1 ;
        RECT 21.424 11.892 21.456 12.636 ;
  LAYER M1 ;
        RECT 21.424 12.732 21.456 12.972 ;
  LAYER M1 ;
        RECT 21.424 13.068 21.456 13.812 ;
  LAYER M1 ;
        RECT 21.424 13.908 21.456 14.148 ;
  LAYER M1 ;
        RECT 21.424 14.244 21.456 14.988 ;
  LAYER M1 ;
        RECT 21.424 15.084 21.456 15.324 ;
  LAYER M1 ;
        RECT 21.424 15.42 21.456 16.164 ;
  LAYER M1 ;
        RECT 21.424 16.26 21.456 16.5 ;
  LAYER M1 ;
        RECT 21.424 16.596 21.456 17.34 ;
  LAYER M1 ;
        RECT 21.424 17.436 21.456 17.676 ;
  LAYER M1 ;
        RECT 21.424 17.94 21.456 18.18 ;
  LAYER M1 ;
        RECT 21.344 9.54 21.376 10.284 ;
  LAYER M1 ;
        RECT 21.344 10.716 21.376 11.46 ;
  LAYER M1 ;
        RECT 21.344 11.892 21.376 12.636 ;
  LAYER M1 ;
        RECT 21.344 13.068 21.376 13.812 ;
  LAYER M1 ;
        RECT 21.344 14.244 21.376 14.988 ;
  LAYER M1 ;
        RECT 21.344 15.42 21.376 16.164 ;
  LAYER M1 ;
        RECT 21.344 16.596 21.376 17.34 ;
  LAYER M1 ;
        RECT 21.504 9.54 21.536 10.284 ;
  LAYER M1 ;
        RECT 21.504 10.716 21.536 11.46 ;
  LAYER M1 ;
        RECT 21.504 11.892 21.536 12.636 ;
  LAYER M1 ;
        RECT 21.504 13.068 21.536 13.812 ;
  LAYER M1 ;
        RECT 21.504 14.244 21.536 14.988 ;
  LAYER M1 ;
        RECT 21.504 15.42 21.536 16.164 ;
  LAYER M1 ;
        RECT 21.504 16.596 21.536 17.34 ;
  LAYER M1 ;
        RECT 22.064 9.54 22.096 10.284 ;
  LAYER M1 ;
        RECT 22.064 10.38 22.096 10.62 ;
  LAYER M1 ;
        RECT 22.064 10.716 22.096 11.46 ;
  LAYER M1 ;
        RECT 22.064 11.556 22.096 11.796 ;
  LAYER M1 ;
        RECT 22.064 11.892 22.096 12.636 ;
  LAYER M1 ;
        RECT 22.064 12.732 22.096 12.972 ;
  LAYER M1 ;
        RECT 22.064 13.068 22.096 13.812 ;
  LAYER M1 ;
        RECT 22.064 13.908 22.096 14.148 ;
  LAYER M1 ;
        RECT 22.064 14.244 22.096 14.988 ;
  LAYER M1 ;
        RECT 22.064 15.084 22.096 15.324 ;
  LAYER M1 ;
        RECT 22.064 15.42 22.096 16.164 ;
  LAYER M1 ;
        RECT 22.064 16.26 22.096 16.5 ;
  LAYER M1 ;
        RECT 22.064 16.596 22.096 17.34 ;
  LAYER M1 ;
        RECT 22.064 17.436 22.096 17.676 ;
  LAYER M1 ;
        RECT 22.064 17.94 22.096 18.18 ;
  LAYER M1 ;
        RECT 21.984 9.54 22.016 10.284 ;
  LAYER M1 ;
        RECT 21.984 10.716 22.016 11.46 ;
  LAYER M1 ;
        RECT 21.984 11.892 22.016 12.636 ;
  LAYER M1 ;
        RECT 21.984 13.068 22.016 13.812 ;
  LAYER M1 ;
        RECT 21.984 14.244 22.016 14.988 ;
  LAYER M1 ;
        RECT 21.984 15.42 22.016 16.164 ;
  LAYER M1 ;
        RECT 21.984 16.596 22.016 17.34 ;
  LAYER M1 ;
        RECT 22.144 9.54 22.176 10.284 ;
  LAYER M1 ;
        RECT 22.144 10.716 22.176 11.46 ;
  LAYER M1 ;
        RECT 22.144 11.892 22.176 12.636 ;
  LAYER M1 ;
        RECT 22.144 13.068 22.176 13.812 ;
  LAYER M1 ;
        RECT 22.144 14.244 22.176 14.988 ;
  LAYER M1 ;
        RECT 22.144 15.42 22.176 16.164 ;
  LAYER M1 ;
        RECT 22.144 16.596 22.176 17.34 ;
  LAYER M1 ;
        RECT 22.704 9.54 22.736 10.284 ;
  LAYER M1 ;
        RECT 22.704 10.38 22.736 10.62 ;
  LAYER M1 ;
        RECT 22.704 10.716 22.736 11.46 ;
  LAYER M1 ;
        RECT 22.704 11.556 22.736 11.796 ;
  LAYER M1 ;
        RECT 22.704 11.892 22.736 12.636 ;
  LAYER M1 ;
        RECT 22.704 12.732 22.736 12.972 ;
  LAYER M1 ;
        RECT 22.704 13.068 22.736 13.812 ;
  LAYER M1 ;
        RECT 22.704 13.908 22.736 14.148 ;
  LAYER M1 ;
        RECT 22.704 14.244 22.736 14.988 ;
  LAYER M1 ;
        RECT 22.704 15.084 22.736 15.324 ;
  LAYER M1 ;
        RECT 22.704 15.42 22.736 16.164 ;
  LAYER M1 ;
        RECT 22.704 16.26 22.736 16.5 ;
  LAYER M1 ;
        RECT 22.704 16.596 22.736 17.34 ;
  LAYER M1 ;
        RECT 22.704 17.436 22.736 17.676 ;
  LAYER M1 ;
        RECT 22.704 17.94 22.736 18.18 ;
  LAYER M1 ;
        RECT 22.624 9.54 22.656 10.284 ;
  LAYER M1 ;
        RECT 22.624 10.716 22.656 11.46 ;
  LAYER M1 ;
        RECT 22.624 11.892 22.656 12.636 ;
  LAYER M1 ;
        RECT 22.624 13.068 22.656 13.812 ;
  LAYER M1 ;
        RECT 22.624 14.244 22.656 14.988 ;
  LAYER M1 ;
        RECT 22.624 15.42 22.656 16.164 ;
  LAYER M1 ;
        RECT 22.624 16.596 22.656 17.34 ;
  LAYER M1 ;
        RECT 22.784 9.54 22.816 10.284 ;
  LAYER M1 ;
        RECT 22.784 10.716 22.816 11.46 ;
  LAYER M1 ;
        RECT 22.784 11.892 22.816 12.636 ;
  LAYER M1 ;
        RECT 22.784 13.068 22.816 13.812 ;
  LAYER M1 ;
        RECT 22.784 14.244 22.816 14.988 ;
  LAYER M1 ;
        RECT 22.784 15.42 22.816 16.164 ;
  LAYER M1 ;
        RECT 22.784 16.596 22.816 17.34 ;
  LAYER M1 ;
        RECT 23.344 9.54 23.376 10.284 ;
  LAYER M1 ;
        RECT 23.344 10.38 23.376 10.62 ;
  LAYER M1 ;
        RECT 23.344 10.716 23.376 11.46 ;
  LAYER M1 ;
        RECT 23.344 11.556 23.376 11.796 ;
  LAYER M1 ;
        RECT 23.344 11.892 23.376 12.636 ;
  LAYER M1 ;
        RECT 23.344 12.732 23.376 12.972 ;
  LAYER M1 ;
        RECT 23.344 13.068 23.376 13.812 ;
  LAYER M1 ;
        RECT 23.344 13.908 23.376 14.148 ;
  LAYER M1 ;
        RECT 23.344 14.244 23.376 14.988 ;
  LAYER M1 ;
        RECT 23.344 15.084 23.376 15.324 ;
  LAYER M1 ;
        RECT 23.344 15.42 23.376 16.164 ;
  LAYER M1 ;
        RECT 23.344 16.26 23.376 16.5 ;
  LAYER M1 ;
        RECT 23.344 16.596 23.376 17.34 ;
  LAYER M1 ;
        RECT 23.344 17.436 23.376 17.676 ;
  LAYER M1 ;
        RECT 23.344 17.94 23.376 18.18 ;
  LAYER M1 ;
        RECT 23.264 9.54 23.296 10.284 ;
  LAYER M1 ;
        RECT 23.264 10.716 23.296 11.46 ;
  LAYER M1 ;
        RECT 23.264 11.892 23.296 12.636 ;
  LAYER M1 ;
        RECT 23.264 13.068 23.296 13.812 ;
  LAYER M1 ;
        RECT 23.264 14.244 23.296 14.988 ;
  LAYER M1 ;
        RECT 23.264 15.42 23.296 16.164 ;
  LAYER M1 ;
        RECT 23.264 16.596 23.296 17.34 ;
  LAYER M1 ;
        RECT 23.424 9.54 23.456 10.284 ;
  LAYER M1 ;
        RECT 23.424 10.716 23.456 11.46 ;
  LAYER M1 ;
        RECT 23.424 11.892 23.456 12.636 ;
  LAYER M1 ;
        RECT 23.424 13.068 23.456 13.812 ;
  LAYER M1 ;
        RECT 23.424 14.244 23.456 14.988 ;
  LAYER M1 ;
        RECT 23.424 15.42 23.456 16.164 ;
  LAYER M1 ;
        RECT 23.424 16.596 23.456 17.34 ;
  LAYER M1 ;
        RECT 23.984 9.54 24.016 10.284 ;
  LAYER M1 ;
        RECT 23.984 10.38 24.016 10.62 ;
  LAYER M1 ;
        RECT 23.984 10.716 24.016 11.46 ;
  LAYER M1 ;
        RECT 23.984 11.556 24.016 11.796 ;
  LAYER M1 ;
        RECT 23.984 11.892 24.016 12.636 ;
  LAYER M1 ;
        RECT 23.984 12.732 24.016 12.972 ;
  LAYER M1 ;
        RECT 23.984 13.068 24.016 13.812 ;
  LAYER M1 ;
        RECT 23.984 13.908 24.016 14.148 ;
  LAYER M1 ;
        RECT 23.984 14.244 24.016 14.988 ;
  LAYER M1 ;
        RECT 23.984 15.084 24.016 15.324 ;
  LAYER M1 ;
        RECT 23.984 15.42 24.016 16.164 ;
  LAYER M1 ;
        RECT 23.984 16.26 24.016 16.5 ;
  LAYER M1 ;
        RECT 23.984 16.596 24.016 17.34 ;
  LAYER M1 ;
        RECT 23.984 17.436 24.016 17.676 ;
  LAYER M1 ;
        RECT 23.984 17.94 24.016 18.18 ;
  LAYER M1 ;
        RECT 23.904 9.54 23.936 10.284 ;
  LAYER M1 ;
        RECT 23.904 10.716 23.936 11.46 ;
  LAYER M1 ;
        RECT 23.904 11.892 23.936 12.636 ;
  LAYER M1 ;
        RECT 23.904 13.068 23.936 13.812 ;
  LAYER M1 ;
        RECT 23.904 14.244 23.936 14.988 ;
  LAYER M1 ;
        RECT 23.904 15.42 23.936 16.164 ;
  LAYER M1 ;
        RECT 23.904 16.596 23.936 17.34 ;
  LAYER M1 ;
        RECT 24.064 9.54 24.096 10.284 ;
  LAYER M1 ;
        RECT 24.064 10.716 24.096 11.46 ;
  LAYER M1 ;
        RECT 24.064 11.892 24.096 12.636 ;
  LAYER M1 ;
        RECT 24.064 13.068 24.096 13.812 ;
  LAYER M1 ;
        RECT 24.064 14.244 24.096 14.988 ;
  LAYER M1 ;
        RECT 24.064 15.42 24.096 16.164 ;
  LAYER M1 ;
        RECT 24.064 16.596 24.096 17.34 ;
  LAYER M1 ;
        RECT 24.624 9.54 24.656 10.284 ;
  LAYER M1 ;
        RECT 24.624 10.38 24.656 10.62 ;
  LAYER M1 ;
        RECT 24.624 10.716 24.656 11.46 ;
  LAYER M1 ;
        RECT 24.624 11.556 24.656 11.796 ;
  LAYER M1 ;
        RECT 24.624 11.892 24.656 12.636 ;
  LAYER M1 ;
        RECT 24.624 12.732 24.656 12.972 ;
  LAYER M1 ;
        RECT 24.624 13.068 24.656 13.812 ;
  LAYER M1 ;
        RECT 24.624 13.908 24.656 14.148 ;
  LAYER M1 ;
        RECT 24.624 14.244 24.656 14.988 ;
  LAYER M1 ;
        RECT 24.624 15.084 24.656 15.324 ;
  LAYER M1 ;
        RECT 24.624 15.42 24.656 16.164 ;
  LAYER M1 ;
        RECT 24.624 16.26 24.656 16.5 ;
  LAYER M1 ;
        RECT 24.624 16.596 24.656 17.34 ;
  LAYER M1 ;
        RECT 24.624 17.436 24.656 17.676 ;
  LAYER M1 ;
        RECT 24.624 17.94 24.656 18.18 ;
  LAYER M1 ;
        RECT 24.544 9.54 24.576 10.284 ;
  LAYER M1 ;
        RECT 24.544 10.716 24.576 11.46 ;
  LAYER M1 ;
        RECT 24.544 11.892 24.576 12.636 ;
  LAYER M1 ;
        RECT 24.544 13.068 24.576 13.812 ;
  LAYER M1 ;
        RECT 24.544 14.244 24.576 14.988 ;
  LAYER M1 ;
        RECT 24.544 15.42 24.576 16.164 ;
  LAYER M1 ;
        RECT 24.544 16.596 24.576 17.34 ;
  LAYER M1 ;
        RECT 24.704 9.54 24.736 10.284 ;
  LAYER M1 ;
        RECT 24.704 10.716 24.736 11.46 ;
  LAYER M1 ;
        RECT 24.704 11.892 24.736 12.636 ;
  LAYER M1 ;
        RECT 24.704 13.068 24.736 13.812 ;
  LAYER M1 ;
        RECT 24.704 14.244 24.736 14.988 ;
  LAYER M1 ;
        RECT 24.704 15.42 24.736 16.164 ;
  LAYER M1 ;
        RECT 24.704 16.596 24.736 17.34 ;
  LAYER M2 ;
        RECT 9.804 9.56 24.756 9.592 ;
  LAYER M2 ;
        RECT 10.444 9.644 24.116 9.676 ;
  LAYER M2 ;
        RECT 9.884 9.728 24.676 9.76 ;
  LAYER M2 ;
        RECT 9.884 10.4 24.676 10.432 ;
  LAYER M2 ;
        RECT 10.524 9.812 24.036 9.844 ;
  LAYER M2 ;
        RECT 10.444 10.736 24.116 10.768 ;
  LAYER M2 ;
        RECT 9.804 10.82 24.756 10.852 ;
  LAYER M2 ;
        RECT 10.524 10.904 24.036 10.936 ;
  LAYER M2 ;
        RECT 9.884 11.576 24.676 11.608 ;
  LAYER M2 ;
        RECT 9.884 10.988 24.676 11.02 ;
  LAYER M2 ;
        RECT 9.804 11.912 24.756 11.944 ;
  LAYER M2 ;
        RECT 10.444 11.996 24.116 12.028 ;
  LAYER M2 ;
        RECT 9.884 12.08 24.676 12.112 ;
  LAYER M2 ;
        RECT 9.884 12.752 24.676 12.784 ;
  LAYER M2 ;
        RECT 10.524 12.164 24.036 12.196 ;
  LAYER M2 ;
        RECT 10.444 13.088 24.116 13.12 ;
  LAYER M2 ;
        RECT 9.804 13.172 24.756 13.204 ;
  LAYER M2 ;
        RECT 10.524 13.256 24.036 13.288 ;
  LAYER M2 ;
        RECT 9.884 13.928 24.676 13.96 ;
  LAYER M2 ;
        RECT 9.884 13.34 24.676 13.372 ;
  LAYER M2 ;
        RECT 9.804 14.264 24.756 14.296 ;
  LAYER M2 ;
        RECT 10.444 14.348 24.116 14.38 ;
  LAYER M2 ;
        RECT 9.884 14.432 24.676 14.464 ;
  LAYER M2 ;
        RECT 9.884 15.104 24.676 15.136 ;
  LAYER M2 ;
        RECT 10.524 14.516 24.036 14.548 ;
  LAYER M2 ;
        RECT 10.444 15.44 24.116 15.472 ;
  LAYER M2 ;
        RECT 9.804 15.524 24.756 15.556 ;
  LAYER M2 ;
        RECT 10.524 15.608 24.036 15.64 ;
  LAYER M2 ;
        RECT 9.884 16.28 24.676 16.312 ;
  LAYER M2 ;
        RECT 9.884 15.692 24.676 15.724 ;
  LAYER M2 ;
        RECT 9.804 16.616 24.756 16.648 ;
  LAYER M2 ;
        RECT 10.444 16.7 24.116 16.732 ;
  LAYER M2 ;
        RECT 9.884 16.784 24.676 16.816 ;
  LAYER M2 ;
        RECT 9.884 17.456 24.676 17.488 ;
  LAYER M2 ;
        RECT 10.524 16.868 24.036 16.9 ;
  LAYER M1 ;
        RECT 0.384 22.476 0.416 23.22 ;
  LAYER M1 ;
        RECT 0.384 23.316 0.416 23.556 ;
  LAYER M1 ;
        RECT 0.384 23.652 0.416 24.396 ;
  LAYER M1 ;
        RECT 0.384 24.492 0.416 24.732 ;
  LAYER M1 ;
        RECT 0.384 24.828 0.416 25.572 ;
  LAYER M1 ;
        RECT 0.384 25.668 0.416 25.908 ;
  LAYER M1 ;
        RECT 0.384 26.004 0.416 26.748 ;
  LAYER M1 ;
        RECT 0.384 26.844 0.416 27.084 ;
  LAYER M1 ;
        RECT 0.384 27.18 0.416 27.924 ;
  LAYER M1 ;
        RECT 0.384 28.02 0.416 28.26 ;
  LAYER M1 ;
        RECT 0.384 28.356 0.416 29.1 ;
  LAYER M1 ;
        RECT 0.384 29.196 0.416 29.436 ;
  LAYER M1 ;
        RECT 0.384 29.532 0.416 30.276 ;
  LAYER M1 ;
        RECT 0.384 30.372 0.416 30.612 ;
  LAYER M1 ;
        RECT 0.384 30.876 0.416 31.116 ;
  LAYER M1 ;
        RECT 0.304 22.476 0.336 23.22 ;
  LAYER M1 ;
        RECT 0.304 23.652 0.336 24.396 ;
  LAYER M1 ;
        RECT 0.304 24.828 0.336 25.572 ;
  LAYER M1 ;
        RECT 0.304 26.004 0.336 26.748 ;
  LAYER M1 ;
        RECT 0.304 27.18 0.336 27.924 ;
  LAYER M1 ;
        RECT 0.304 28.356 0.336 29.1 ;
  LAYER M1 ;
        RECT 0.304 29.532 0.336 30.276 ;
  LAYER M1 ;
        RECT 0.464 22.476 0.496 23.22 ;
  LAYER M1 ;
        RECT 0.464 23.652 0.496 24.396 ;
  LAYER M1 ;
        RECT 0.464 24.828 0.496 25.572 ;
  LAYER M1 ;
        RECT 0.464 26.004 0.496 26.748 ;
  LAYER M1 ;
        RECT 0.464 27.18 0.496 27.924 ;
  LAYER M1 ;
        RECT 0.464 28.356 0.496 29.1 ;
  LAYER M1 ;
        RECT 0.464 29.532 0.496 30.276 ;
  LAYER M1 ;
        RECT 1.024 22.476 1.056 23.22 ;
  LAYER M1 ;
        RECT 1.024 23.316 1.056 23.556 ;
  LAYER M1 ;
        RECT 1.024 23.652 1.056 24.396 ;
  LAYER M1 ;
        RECT 1.024 24.492 1.056 24.732 ;
  LAYER M1 ;
        RECT 1.024 24.828 1.056 25.572 ;
  LAYER M1 ;
        RECT 1.024 25.668 1.056 25.908 ;
  LAYER M1 ;
        RECT 1.024 26.004 1.056 26.748 ;
  LAYER M1 ;
        RECT 1.024 26.844 1.056 27.084 ;
  LAYER M1 ;
        RECT 1.024 27.18 1.056 27.924 ;
  LAYER M1 ;
        RECT 1.024 28.02 1.056 28.26 ;
  LAYER M1 ;
        RECT 1.024 28.356 1.056 29.1 ;
  LAYER M1 ;
        RECT 1.024 29.196 1.056 29.436 ;
  LAYER M1 ;
        RECT 1.024 29.532 1.056 30.276 ;
  LAYER M1 ;
        RECT 1.024 30.372 1.056 30.612 ;
  LAYER M1 ;
        RECT 1.024 30.876 1.056 31.116 ;
  LAYER M1 ;
        RECT 0.944 22.476 0.976 23.22 ;
  LAYER M1 ;
        RECT 0.944 23.652 0.976 24.396 ;
  LAYER M1 ;
        RECT 0.944 24.828 0.976 25.572 ;
  LAYER M1 ;
        RECT 0.944 26.004 0.976 26.748 ;
  LAYER M1 ;
        RECT 0.944 27.18 0.976 27.924 ;
  LAYER M1 ;
        RECT 0.944 28.356 0.976 29.1 ;
  LAYER M1 ;
        RECT 0.944 29.532 0.976 30.276 ;
  LAYER M1 ;
        RECT 1.104 22.476 1.136 23.22 ;
  LAYER M1 ;
        RECT 1.104 23.652 1.136 24.396 ;
  LAYER M1 ;
        RECT 1.104 24.828 1.136 25.572 ;
  LAYER M1 ;
        RECT 1.104 26.004 1.136 26.748 ;
  LAYER M1 ;
        RECT 1.104 27.18 1.136 27.924 ;
  LAYER M1 ;
        RECT 1.104 28.356 1.136 29.1 ;
  LAYER M1 ;
        RECT 1.104 29.532 1.136 30.276 ;
  LAYER M1 ;
        RECT 1.664 22.476 1.696 23.22 ;
  LAYER M1 ;
        RECT 1.664 23.316 1.696 23.556 ;
  LAYER M1 ;
        RECT 1.664 23.652 1.696 24.396 ;
  LAYER M1 ;
        RECT 1.664 24.492 1.696 24.732 ;
  LAYER M1 ;
        RECT 1.664 24.828 1.696 25.572 ;
  LAYER M1 ;
        RECT 1.664 25.668 1.696 25.908 ;
  LAYER M1 ;
        RECT 1.664 26.004 1.696 26.748 ;
  LAYER M1 ;
        RECT 1.664 26.844 1.696 27.084 ;
  LAYER M1 ;
        RECT 1.664 27.18 1.696 27.924 ;
  LAYER M1 ;
        RECT 1.664 28.02 1.696 28.26 ;
  LAYER M1 ;
        RECT 1.664 28.356 1.696 29.1 ;
  LAYER M1 ;
        RECT 1.664 29.196 1.696 29.436 ;
  LAYER M1 ;
        RECT 1.664 29.532 1.696 30.276 ;
  LAYER M1 ;
        RECT 1.664 30.372 1.696 30.612 ;
  LAYER M1 ;
        RECT 1.664 30.876 1.696 31.116 ;
  LAYER M1 ;
        RECT 1.584 22.476 1.616 23.22 ;
  LAYER M1 ;
        RECT 1.584 23.652 1.616 24.396 ;
  LAYER M1 ;
        RECT 1.584 24.828 1.616 25.572 ;
  LAYER M1 ;
        RECT 1.584 26.004 1.616 26.748 ;
  LAYER M1 ;
        RECT 1.584 27.18 1.616 27.924 ;
  LAYER M1 ;
        RECT 1.584 28.356 1.616 29.1 ;
  LAYER M1 ;
        RECT 1.584 29.532 1.616 30.276 ;
  LAYER M1 ;
        RECT 1.744 22.476 1.776 23.22 ;
  LAYER M1 ;
        RECT 1.744 23.652 1.776 24.396 ;
  LAYER M1 ;
        RECT 1.744 24.828 1.776 25.572 ;
  LAYER M1 ;
        RECT 1.744 26.004 1.776 26.748 ;
  LAYER M1 ;
        RECT 1.744 27.18 1.776 27.924 ;
  LAYER M1 ;
        RECT 1.744 28.356 1.776 29.1 ;
  LAYER M1 ;
        RECT 1.744 29.532 1.776 30.276 ;
  LAYER M1 ;
        RECT 2.304 22.476 2.336 23.22 ;
  LAYER M1 ;
        RECT 2.304 23.316 2.336 23.556 ;
  LAYER M1 ;
        RECT 2.304 23.652 2.336 24.396 ;
  LAYER M1 ;
        RECT 2.304 24.492 2.336 24.732 ;
  LAYER M1 ;
        RECT 2.304 24.828 2.336 25.572 ;
  LAYER M1 ;
        RECT 2.304 25.668 2.336 25.908 ;
  LAYER M1 ;
        RECT 2.304 26.004 2.336 26.748 ;
  LAYER M1 ;
        RECT 2.304 26.844 2.336 27.084 ;
  LAYER M1 ;
        RECT 2.304 27.18 2.336 27.924 ;
  LAYER M1 ;
        RECT 2.304 28.02 2.336 28.26 ;
  LAYER M1 ;
        RECT 2.304 28.356 2.336 29.1 ;
  LAYER M1 ;
        RECT 2.304 29.196 2.336 29.436 ;
  LAYER M1 ;
        RECT 2.304 29.532 2.336 30.276 ;
  LAYER M1 ;
        RECT 2.304 30.372 2.336 30.612 ;
  LAYER M1 ;
        RECT 2.304 30.876 2.336 31.116 ;
  LAYER M1 ;
        RECT 2.224 22.476 2.256 23.22 ;
  LAYER M1 ;
        RECT 2.224 23.652 2.256 24.396 ;
  LAYER M1 ;
        RECT 2.224 24.828 2.256 25.572 ;
  LAYER M1 ;
        RECT 2.224 26.004 2.256 26.748 ;
  LAYER M1 ;
        RECT 2.224 27.18 2.256 27.924 ;
  LAYER M1 ;
        RECT 2.224 28.356 2.256 29.1 ;
  LAYER M1 ;
        RECT 2.224 29.532 2.256 30.276 ;
  LAYER M1 ;
        RECT 2.384 22.476 2.416 23.22 ;
  LAYER M1 ;
        RECT 2.384 23.652 2.416 24.396 ;
  LAYER M1 ;
        RECT 2.384 24.828 2.416 25.572 ;
  LAYER M1 ;
        RECT 2.384 26.004 2.416 26.748 ;
  LAYER M1 ;
        RECT 2.384 27.18 2.416 27.924 ;
  LAYER M1 ;
        RECT 2.384 28.356 2.416 29.1 ;
  LAYER M1 ;
        RECT 2.384 29.532 2.416 30.276 ;
  LAYER M1 ;
        RECT 2.944 22.476 2.976 23.22 ;
  LAYER M1 ;
        RECT 2.944 23.316 2.976 23.556 ;
  LAYER M1 ;
        RECT 2.944 23.652 2.976 24.396 ;
  LAYER M1 ;
        RECT 2.944 24.492 2.976 24.732 ;
  LAYER M1 ;
        RECT 2.944 24.828 2.976 25.572 ;
  LAYER M1 ;
        RECT 2.944 25.668 2.976 25.908 ;
  LAYER M1 ;
        RECT 2.944 26.004 2.976 26.748 ;
  LAYER M1 ;
        RECT 2.944 26.844 2.976 27.084 ;
  LAYER M1 ;
        RECT 2.944 27.18 2.976 27.924 ;
  LAYER M1 ;
        RECT 2.944 28.02 2.976 28.26 ;
  LAYER M1 ;
        RECT 2.944 28.356 2.976 29.1 ;
  LAYER M1 ;
        RECT 2.944 29.196 2.976 29.436 ;
  LAYER M1 ;
        RECT 2.944 29.532 2.976 30.276 ;
  LAYER M1 ;
        RECT 2.944 30.372 2.976 30.612 ;
  LAYER M1 ;
        RECT 2.944 30.876 2.976 31.116 ;
  LAYER M1 ;
        RECT 2.864 22.476 2.896 23.22 ;
  LAYER M1 ;
        RECT 2.864 23.652 2.896 24.396 ;
  LAYER M1 ;
        RECT 2.864 24.828 2.896 25.572 ;
  LAYER M1 ;
        RECT 2.864 26.004 2.896 26.748 ;
  LAYER M1 ;
        RECT 2.864 27.18 2.896 27.924 ;
  LAYER M1 ;
        RECT 2.864 28.356 2.896 29.1 ;
  LAYER M1 ;
        RECT 2.864 29.532 2.896 30.276 ;
  LAYER M1 ;
        RECT 3.024 22.476 3.056 23.22 ;
  LAYER M1 ;
        RECT 3.024 23.652 3.056 24.396 ;
  LAYER M1 ;
        RECT 3.024 24.828 3.056 25.572 ;
  LAYER M1 ;
        RECT 3.024 26.004 3.056 26.748 ;
  LAYER M1 ;
        RECT 3.024 27.18 3.056 27.924 ;
  LAYER M1 ;
        RECT 3.024 28.356 3.056 29.1 ;
  LAYER M1 ;
        RECT 3.024 29.532 3.056 30.276 ;
  LAYER M1 ;
        RECT 3.584 22.476 3.616 23.22 ;
  LAYER M1 ;
        RECT 3.584 23.316 3.616 23.556 ;
  LAYER M1 ;
        RECT 3.584 23.652 3.616 24.396 ;
  LAYER M1 ;
        RECT 3.584 24.492 3.616 24.732 ;
  LAYER M1 ;
        RECT 3.584 24.828 3.616 25.572 ;
  LAYER M1 ;
        RECT 3.584 25.668 3.616 25.908 ;
  LAYER M1 ;
        RECT 3.584 26.004 3.616 26.748 ;
  LAYER M1 ;
        RECT 3.584 26.844 3.616 27.084 ;
  LAYER M1 ;
        RECT 3.584 27.18 3.616 27.924 ;
  LAYER M1 ;
        RECT 3.584 28.02 3.616 28.26 ;
  LAYER M1 ;
        RECT 3.584 28.356 3.616 29.1 ;
  LAYER M1 ;
        RECT 3.584 29.196 3.616 29.436 ;
  LAYER M1 ;
        RECT 3.584 29.532 3.616 30.276 ;
  LAYER M1 ;
        RECT 3.584 30.372 3.616 30.612 ;
  LAYER M1 ;
        RECT 3.584 30.876 3.616 31.116 ;
  LAYER M1 ;
        RECT 3.504 22.476 3.536 23.22 ;
  LAYER M1 ;
        RECT 3.504 23.652 3.536 24.396 ;
  LAYER M1 ;
        RECT 3.504 24.828 3.536 25.572 ;
  LAYER M1 ;
        RECT 3.504 26.004 3.536 26.748 ;
  LAYER M1 ;
        RECT 3.504 27.18 3.536 27.924 ;
  LAYER M1 ;
        RECT 3.504 28.356 3.536 29.1 ;
  LAYER M1 ;
        RECT 3.504 29.532 3.536 30.276 ;
  LAYER M1 ;
        RECT 3.664 22.476 3.696 23.22 ;
  LAYER M1 ;
        RECT 3.664 23.652 3.696 24.396 ;
  LAYER M1 ;
        RECT 3.664 24.828 3.696 25.572 ;
  LAYER M1 ;
        RECT 3.664 26.004 3.696 26.748 ;
  LAYER M1 ;
        RECT 3.664 27.18 3.696 27.924 ;
  LAYER M1 ;
        RECT 3.664 28.356 3.696 29.1 ;
  LAYER M1 ;
        RECT 3.664 29.532 3.696 30.276 ;
  LAYER M1 ;
        RECT 4.224 22.476 4.256 23.22 ;
  LAYER M1 ;
        RECT 4.224 23.316 4.256 23.556 ;
  LAYER M1 ;
        RECT 4.224 23.652 4.256 24.396 ;
  LAYER M1 ;
        RECT 4.224 24.492 4.256 24.732 ;
  LAYER M1 ;
        RECT 4.224 24.828 4.256 25.572 ;
  LAYER M1 ;
        RECT 4.224 25.668 4.256 25.908 ;
  LAYER M1 ;
        RECT 4.224 26.004 4.256 26.748 ;
  LAYER M1 ;
        RECT 4.224 26.844 4.256 27.084 ;
  LAYER M1 ;
        RECT 4.224 27.18 4.256 27.924 ;
  LAYER M1 ;
        RECT 4.224 28.02 4.256 28.26 ;
  LAYER M1 ;
        RECT 4.224 28.356 4.256 29.1 ;
  LAYER M1 ;
        RECT 4.224 29.196 4.256 29.436 ;
  LAYER M1 ;
        RECT 4.224 29.532 4.256 30.276 ;
  LAYER M1 ;
        RECT 4.224 30.372 4.256 30.612 ;
  LAYER M1 ;
        RECT 4.224 30.876 4.256 31.116 ;
  LAYER M1 ;
        RECT 4.144 22.476 4.176 23.22 ;
  LAYER M1 ;
        RECT 4.144 23.652 4.176 24.396 ;
  LAYER M1 ;
        RECT 4.144 24.828 4.176 25.572 ;
  LAYER M1 ;
        RECT 4.144 26.004 4.176 26.748 ;
  LAYER M1 ;
        RECT 4.144 27.18 4.176 27.924 ;
  LAYER M1 ;
        RECT 4.144 28.356 4.176 29.1 ;
  LAYER M1 ;
        RECT 4.144 29.532 4.176 30.276 ;
  LAYER M1 ;
        RECT 4.304 22.476 4.336 23.22 ;
  LAYER M1 ;
        RECT 4.304 23.652 4.336 24.396 ;
  LAYER M1 ;
        RECT 4.304 24.828 4.336 25.572 ;
  LAYER M1 ;
        RECT 4.304 26.004 4.336 26.748 ;
  LAYER M1 ;
        RECT 4.304 27.18 4.336 27.924 ;
  LAYER M1 ;
        RECT 4.304 28.356 4.336 29.1 ;
  LAYER M1 ;
        RECT 4.304 29.532 4.336 30.276 ;
  LAYER M1 ;
        RECT 4.864 22.476 4.896 23.22 ;
  LAYER M1 ;
        RECT 4.864 23.316 4.896 23.556 ;
  LAYER M1 ;
        RECT 4.864 23.652 4.896 24.396 ;
  LAYER M1 ;
        RECT 4.864 24.492 4.896 24.732 ;
  LAYER M1 ;
        RECT 4.864 24.828 4.896 25.572 ;
  LAYER M1 ;
        RECT 4.864 25.668 4.896 25.908 ;
  LAYER M1 ;
        RECT 4.864 26.004 4.896 26.748 ;
  LAYER M1 ;
        RECT 4.864 26.844 4.896 27.084 ;
  LAYER M1 ;
        RECT 4.864 27.18 4.896 27.924 ;
  LAYER M1 ;
        RECT 4.864 28.02 4.896 28.26 ;
  LAYER M1 ;
        RECT 4.864 28.356 4.896 29.1 ;
  LAYER M1 ;
        RECT 4.864 29.196 4.896 29.436 ;
  LAYER M1 ;
        RECT 4.864 29.532 4.896 30.276 ;
  LAYER M1 ;
        RECT 4.864 30.372 4.896 30.612 ;
  LAYER M1 ;
        RECT 4.864 30.876 4.896 31.116 ;
  LAYER M1 ;
        RECT 4.784 22.476 4.816 23.22 ;
  LAYER M1 ;
        RECT 4.784 23.652 4.816 24.396 ;
  LAYER M1 ;
        RECT 4.784 24.828 4.816 25.572 ;
  LAYER M1 ;
        RECT 4.784 26.004 4.816 26.748 ;
  LAYER M1 ;
        RECT 4.784 27.18 4.816 27.924 ;
  LAYER M1 ;
        RECT 4.784 28.356 4.816 29.1 ;
  LAYER M1 ;
        RECT 4.784 29.532 4.816 30.276 ;
  LAYER M1 ;
        RECT 4.944 22.476 4.976 23.22 ;
  LAYER M1 ;
        RECT 4.944 23.652 4.976 24.396 ;
  LAYER M1 ;
        RECT 4.944 24.828 4.976 25.572 ;
  LAYER M1 ;
        RECT 4.944 26.004 4.976 26.748 ;
  LAYER M1 ;
        RECT 4.944 27.18 4.976 27.924 ;
  LAYER M1 ;
        RECT 4.944 28.356 4.976 29.1 ;
  LAYER M1 ;
        RECT 4.944 29.532 4.976 30.276 ;
  LAYER M1 ;
        RECT 5.504 22.476 5.536 23.22 ;
  LAYER M1 ;
        RECT 5.504 23.316 5.536 23.556 ;
  LAYER M1 ;
        RECT 5.504 23.652 5.536 24.396 ;
  LAYER M1 ;
        RECT 5.504 24.492 5.536 24.732 ;
  LAYER M1 ;
        RECT 5.504 24.828 5.536 25.572 ;
  LAYER M1 ;
        RECT 5.504 25.668 5.536 25.908 ;
  LAYER M1 ;
        RECT 5.504 26.004 5.536 26.748 ;
  LAYER M1 ;
        RECT 5.504 26.844 5.536 27.084 ;
  LAYER M1 ;
        RECT 5.504 27.18 5.536 27.924 ;
  LAYER M1 ;
        RECT 5.504 28.02 5.536 28.26 ;
  LAYER M1 ;
        RECT 5.504 28.356 5.536 29.1 ;
  LAYER M1 ;
        RECT 5.504 29.196 5.536 29.436 ;
  LAYER M1 ;
        RECT 5.504 29.532 5.536 30.276 ;
  LAYER M1 ;
        RECT 5.504 30.372 5.536 30.612 ;
  LAYER M1 ;
        RECT 5.504 30.876 5.536 31.116 ;
  LAYER M1 ;
        RECT 5.424 22.476 5.456 23.22 ;
  LAYER M1 ;
        RECT 5.424 23.652 5.456 24.396 ;
  LAYER M1 ;
        RECT 5.424 24.828 5.456 25.572 ;
  LAYER M1 ;
        RECT 5.424 26.004 5.456 26.748 ;
  LAYER M1 ;
        RECT 5.424 27.18 5.456 27.924 ;
  LAYER M1 ;
        RECT 5.424 28.356 5.456 29.1 ;
  LAYER M1 ;
        RECT 5.424 29.532 5.456 30.276 ;
  LAYER M1 ;
        RECT 5.584 22.476 5.616 23.22 ;
  LAYER M1 ;
        RECT 5.584 23.652 5.616 24.396 ;
  LAYER M1 ;
        RECT 5.584 24.828 5.616 25.572 ;
  LAYER M1 ;
        RECT 5.584 26.004 5.616 26.748 ;
  LAYER M1 ;
        RECT 5.584 27.18 5.616 27.924 ;
  LAYER M1 ;
        RECT 5.584 28.356 5.616 29.1 ;
  LAYER M1 ;
        RECT 5.584 29.532 5.616 30.276 ;
  LAYER M1 ;
        RECT 6.144 22.476 6.176 23.22 ;
  LAYER M1 ;
        RECT 6.144 23.316 6.176 23.556 ;
  LAYER M1 ;
        RECT 6.144 23.652 6.176 24.396 ;
  LAYER M1 ;
        RECT 6.144 24.492 6.176 24.732 ;
  LAYER M1 ;
        RECT 6.144 24.828 6.176 25.572 ;
  LAYER M1 ;
        RECT 6.144 25.668 6.176 25.908 ;
  LAYER M1 ;
        RECT 6.144 26.004 6.176 26.748 ;
  LAYER M1 ;
        RECT 6.144 26.844 6.176 27.084 ;
  LAYER M1 ;
        RECT 6.144 27.18 6.176 27.924 ;
  LAYER M1 ;
        RECT 6.144 28.02 6.176 28.26 ;
  LAYER M1 ;
        RECT 6.144 28.356 6.176 29.1 ;
  LAYER M1 ;
        RECT 6.144 29.196 6.176 29.436 ;
  LAYER M1 ;
        RECT 6.144 29.532 6.176 30.276 ;
  LAYER M1 ;
        RECT 6.144 30.372 6.176 30.612 ;
  LAYER M1 ;
        RECT 6.144 30.876 6.176 31.116 ;
  LAYER M1 ;
        RECT 6.064 22.476 6.096 23.22 ;
  LAYER M1 ;
        RECT 6.064 23.652 6.096 24.396 ;
  LAYER M1 ;
        RECT 6.064 24.828 6.096 25.572 ;
  LAYER M1 ;
        RECT 6.064 26.004 6.096 26.748 ;
  LAYER M1 ;
        RECT 6.064 27.18 6.096 27.924 ;
  LAYER M1 ;
        RECT 6.064 28.356 6.096 29.1 ;
  LAYER M1 ;
        RECT 6.064 29.532 6.096 30.276 ;
  LAYER M1 ;
        RECT 6.224 22.476 6.256 23.22 ;
  LAYER M1 ;
        RECT 6.224 23.652 6.256 24.396 ;
  LAYER M1 ;
        RECT 6.224 24.828 6.256 25.572 ;
  LAYER M1 ;
        RECT 6.224 26.004 6.256 26.748 ;
  LAYER M1 ;
        RECT 6.224 27.18 6.256 27.924 ;
  LAYER M1 ;
        RECT 6.224 28.356 6.256 29.1 ;
  LAYER M1 ;
        RECT 6.224 29.532 6.256 30.276 ;
  LAYER M1 ;
        RECT 6.784 22.476 6.816 23.22 ;
  LAYER M1 ;
        RECT 6.784 23.316 6.816 23.556 ;
  LAYER M1 ;
        RECT 6.784 23.652 6.816 24.396 ;
  LAYER M1 ;
        RECT 6.784 24.492 6.816 24.732 ;
  LAYER M1 ;
        RECT 6.784 24.828 6.816 25.572 ;
  LAYER M1 ;
        RECT 6.784 25.668 6.816 25.908 ;
  LAYER M1 ;
        RECT 6.784 26.004 6.816 26.748 ;
  LAYER M1 ;
        RECT 6.784 26.844 6.816 27.084 ;
  LAYER M1 ;
        RECT 6.784 27.18 6.816 27.924 ;
  LAYER M1 ;
        RECT 6.784 28.02 6.816 28.26 ;
  LAYER M1 ;
        RECT 6.784 28.356 6.816 29.1 ;
  LAYER M1 ;
        RECT 6.784 29.196 6.816 29.436 ;
  LAYER M1 ;
        RECT 6.784 29.532 6.816 30.276 ;
  LAYER M1 ;
        RECT 6.784 30.372 6.816 30.612 ;
  LAYER M1 ;
        RECT 6.784 30.876 6.816 31.116 ;
  LAYER M1 ;
        RECT 6.704 22.476 6.736 23.22 ;
  LAYER M1 ;
        RECT 6.704 23.652 6.736 24.396 ;
  LAYER M1 ;
        RECT 6.704 24.828 6.736 25.572 ;
  LAYER M1 ;
        RECT 6.704 26.004 6.736 26.748 ;
  LAYER M1 ;
        RECT 6.704 27.18 6.736 27.924 ;
  LAYER M1 ;
        RECT 6.704 28.356 6.736 29.1 ;
  LAYER M1 ;
        RECT 6.704 29.532 6.736 30.276 ;
  LAYER M1 ;
        RECT 6.864 22.476 6.896 23.22 ;
  LAYER M1 ;
        RECT 6.864 23.652 6.896 24.396 ;
  LAYER M1 ;
        RECT 6.864 24.828 6.896 25.572 ;
  LAYER M1 ;
        RECT 6.864 26.004 6.896 26.748 ;
  LAYER M1 ;
        RECT 6.864 27.18 6.896 27.924 ;
  LAYER M1 ;
        RECT 6.864 28.356 6.896 29.1 ;
  LAYER M1 ;
        RECT 6.864 29.532 6.896 30.276 ;
  LAYER M1 ;
        RECT 7.424 22.476 7.456 23.22 ;
  LAYER M1 ;
        RECT 7.424 23.316 7.456 23.556 ;
  LAYER M1 ;
        RECT 7.424 23.652 7.456 24.396 ;
  LAYER M1 ;
        RECT 7.424 24.492 7.456 24.732 ;
  LAYER M1 ;
        RECT 7.424 24.828 7.456 25.572 ;
  LAYER M1 ;
        RECT 7.424 25.668 7.456 25.908 ;
  LAYER M1 ;
        RECT 7.424 26.004 7.456 26.748 ;
  LAYER M1 ;
        RECT 7.424 26.844 7.456 27.084 ;
  LAYER M1 ;
        RECT 7.424 27.18 7.456 27.924 ;
  LAYER M1 ;
        RECT 7.424 28.02 7.456 28.26 ;
  LAYER M1 ;
        RECT 7.424 28.356 7.456 29.1 ;
  LAYER M1 ;
        RECT 7.424 29.196 7.456 29.436 ;
  LAYER M1 ;
        RECT 7.424 29.532 7.456 30.276 ;
  LAYER M1 ;
        RECT 7.424 30.372 7.456 30.612 ;
  LAYER M1 ;
        RECT 7.424 30.876 7.456 31.116 ;
  LAYER M1 ;
        RECT 7.344 22.476 7.376 23.22 ;
  LAYER M1 ;
        RECT 7.344 23.652 7.376 24.396 ;
  LAYER M1 ;
        RECT 7.344 24.828 7.376 25.572 ;
  LAYER M1 ;
        RECT 7.344 26.004 7.376 26.748 ;
  LAYER M1 ;
        RECT 7.344 27.18 7.376 27.924 ;
  LAYER M1 ;
        RECT 7.344 28.356 7.376 29.1 ;
  LAYER M1 ;
        RECT 7.344 29.532 7.376 30.276 ;
  LAYER M1 ;
        RECT 7.504 22.476 7.536 23.22 ;
  LAYER M1 ;
        RECT 7.504 23.652 7.536 24.396 ;
  LAYER M1 ;
        RECT 7.504 24.828 7.536 25.572 ;
  LAYER M1 ;
        RECT 7.504 26.004 7.536 26.748 ;
  LAYER M1 ;
        RECT 7.504 27.18 7.536 27.924 ;
  LAYER M1 ;
        RECT 7.504 28.356 7.536 29.1 ;
  LAYER M1 ;
        RECT 7.504 29.532 7.536 30.276 ;
  LAYER M1 ;
        RECT 8.064 22.476 8.096 23.22 ;
  LAYER M1 ;
        RECT 8.064 23.316 8.096 23.556 ;
  LAYER M1 ;
        RECT 8.064 23.652 8.096 24.396 ;
  LAYER M1 ;
        RECT 8.064 24.492 8.096 24.732 ;
  LAYER M1 ;
        RECT 8.064 24.828 8.096 25.572 ;
  LAYER M1 ;
        RECT 8.064 25.668 8.096 25.908 ;
  LAYER M1 ;
        RECT 8.064 26.004 8.096 26.748 ;
  LAYER M1 ;
        RECT 8.064 26.844 8.096 27.084 ;
  LAYER M1 ;
        RECT 8.064 27.18 8.096 27.924 ;
  LAYER M1 ;
        RECT 8.064 28.02 8.096 28.26 ;
  LAYER M1 ;
        RECT 8.064 28.356 8.096 29.1 ;
  LAYER M1 ;
        RECT 8.064 29.196 8.096 29.436 ;
  LAYER M1 ;
        RECT 8.064 29.532 8.096 30.276 ;
  LAYER M1 ;
        RECT 8.064 30.372 8.096 30.612 ;
  LAYER M1 ;
        RECT 8.064 30.876 8.096 31.116 ;
  LAYER M1 ;
        RECT 7.984 22.476 8.016 23.22 ;
  LAYER M1 ;
        RECT 7.984 23.652 8.016 24.396 ;
  LAYER M1 ;
        RECT 7.984 24.828 8.016 25.572 ;
  LAYER M1 ;
        RECT 7.984 26.004 8.016 26.748 ;
  LAYER M1 ;
        RECT 7.984 27.18 8.016 27.924 ;
  LAYER M1 ;
        RECT 7.984 28.356 8.016 29.1 ;
  LAYER M1 ;
        RECT 7.984 29.532 8.016 30.276 ;
  LAYER M1 ;
        RECT 8.144 22.476 8.176 23.22 ;
  LAYER M1 ;
        RECT 8.144 23.652 8.176 24.396 ;
  LAYER M1 ;
        RECT 8.144 24.828 8.176 25.572 ;
  LAYER M1 ;
        RECT 8.144 26.004 8.176 26.748 ;
  LAYER M1 ;
        RECT 8.144 27.18 8.176 27.924 ;
  LAYER M1 ;
        RECT 8.144 28.356 8.176 29.1 ;
  LAYER M1 ;
        RECT 8.144 29.532 8.176 30.276 ;
  LAYER M1 ;
        RECT 8.704 22.476 8.736 23.22 ;
  LAYER M1 ;
        RECT 8.704 23.316 8.736 23.556 ;
  LAYER M1 ;
        RECT 8.704 23.652 8.736 24.396 ;
  LAYER M1 ;
        RECT 8.704 24.492 8.736 24.732 ;
  LAYER M1 ;
        RECT 8.704 24.828 8.736 25.572 ;
  LAYER M1 ;
        RECT 8.704 25.668 8.736 25.908 ;
  LAYER M1 ;
        RECT 8.704 26.004 8.736 26.748 ;
  LAYER M1 ;
        RECT 8.704 26.844 8.736 27.084 ;
  LAYER M1 ;
        RECT 8.704 27.18 8.736 27.924 ;
  LAYER M1 ;
        RECT 8.704 28.02 8.736 28.26 ;
  LAYER M1 ;
        RECT 8.704 28.356 8.736 29.1 ;
  LAYER M1 ;
        RECT 8.704 29.196 8.736 29.436 ;
  LAYER M1 ;
        RECT 8.704 29.532 8.736 30.276 ;
  LAYER M1 ;
        RECT 8.704 30.372 8.736 30.612 ;
  LAYER M1 ;
        RECT 8.704 30.876 8.736 31.116 ;
  LAYER M1 ;
        RECT 8.624 22.476 8.656 23.22 ;
  LAYER M1 ;
        RECT 8.624 23.652 8.656 24.396 ;
  LAYER M1 ;
        RECT 8.624 24.828 8.656 25.572 ;
  LAYER M1 ;
        RECT 8.624 26.004 8.656 26.748 ;
  LAYER M1 ;
        RECT 8.624 27.18 8.656 27.924 ;
  LAYER M1 ;
        RECT 8.624 28.356 8.656 29.1 ;
  LAYER M1 ;
        RECT 8.624 29.532 8.656 30.276 ;
  LAYER M1 ;
        RECT 8.784 22.476 8.816 23.22 ;
  LAYER M1 ;
        RECT 8.784 23.652 8.816 24.396 ;
  LAYER M1 ;
        RECT 8.784 24.828 8.816 25.572 ;
  LAYER M1 ;
        RECT 8.784 26.004 8.816 26.748 ;
  LAYER M1 ;
        RECT 8.784 27.18 8.816 27.924 ;
  LAYER M1 ;
        RECT 8.784 28.356 8.816 29.1 ;
  LAYER M1 ;
        RECT 8.784 29.532 8.816 30.276 ;
  LAYER M1 ;
        RECT 9.344 22.476 9.376 23.22 ;
  LAYER M1 ;
        RECT 9.344 23.316 9.376 23.556 ;
  LAYER M1 ;
        RECT 9.344 23.652 9.376 24.396 ;
  LAYER M1 ;
        RECT 9.344 24.492 9.376 24.732 ;
  LAYER M1 ;
        RECT 9.344 24.828 9.376 25.572 ;
  LAYER M1 ;
        RECT 9.344 25.668 9.376 25.908 ;
  LAYER M1 ;
        RECT 9.344 26.004 9.376 26.748 ;
  LAYER M1 ;
        RECT 9.344 26.844 9.376 27.084 ;
  LAYER M1 ;
        RECT 9.344 27.18 9.376 27.924 ;
  LAYER M1 ;
        RECT 9.344 28.02 9.376 28.26 ;
  LAYER M1 ;
        RECT 9.344 28.356 9.376 29.1 ;
  LAYER M1 ;
        RECT 9.344 29.196 9.376 29.436 ;
  LAYER M1 ;
        RECT 9.344 29.532 9.376 30.276 ;
  LAYER M1 ;
        RECT 9.344 30.372 9.376 30.612 ;
  LAYER M1 ;
        RECT 9.344 30.876 9.376 31.116 ;
  LAYER M1 ;
        RECT 9.264 22.476 9.296 23.22 ;
  LAYER M1 ;
        RECT 9.264 23.652 9.296 24.396 ;
  LAYER M1 ;
        RECT 9.264 24.828 9.296 25.572 ;
  LAYER M1 ;
        RECT 9.264 26.004 9.296 26.748 ;
  LAYER M1 ;
        RECT 9.264 27.18 9.296 27.924 ;
  LAYER M1 ;
        RECT 9.264 28.356 9.296 29.1 ;
  LAYER M1 ;
        RECT 9.264 29.532 9.296 30.276 ;
  LAYER M1 ;
        RECT 9.424 22.476 9.456 23.22 ;
  LAYER M1 ;
        RECT 9.424 23.652 9.456 24.396 ;
  LAYER M1 ;
        RECT 9.424 24.828 9.456 25.572 ;
  LAYER M1 ;
        RECT 9.424 26.004 9.456 26.748 ;
  LAYER M1 ;
        RECT 9.424 27.18 9.456 27.924 ;
  LAYER M1 ;
        RECT 9.424 28.356 9.456 29.1 ;
  LAYER M1 ;
        RECT 9.424 29.532 9.456 30.276 ;
  LAYER M1 ;
        RECT 9.984 22.476 10.016 23.22 ;
  LAYER M1 ;
        RECT 9.984 23.316 10.016 23.556 ;
  LAYER M1 ;
        RECT 9.984 23.652 10.016 24.396 ;
  LAYER M1 ;
        RECT 9.984 24.492 10.016 24.732 ;
  LAYER M1 ;
        RECT 9.984 24.828 10.016 25.572 ;
  LAYER M1 ;
        RECT 9.984 25.668 10.016 25.908 ;
  LAYER M1 ;
        RECT 9.984 26.004 10.016 26.748 ;
  LAYER M1 ;
        RECT 9.984 26.844 10.016 27.084 ;
  LAYER M1 ;
        RECT 9.984 27.18 10.016 27.924 ;
  LAYER M1 ;
        RECT 9.984 28.02 10.016 28.26 ;
  LAYER M1 ;
        RECT 9.984 28.356 10.016 29.1 ;
  LAYER M1 ;
        RECT 9.984 29.196 10.016 29.436 ;
  LAYER M1 ;
        RECT 9.984 29.532 10.016 30.276 ;
  LAYER M1 ;
        RECT 9.984 30.372 10.016 30.612 ;
  LAYER M1 ;
        RECT 9.984 30.876 10.016 31.116 ;
  LAYER M1 ;
        RECT 9.904 22.476 9.936 23.22 ;
  LAYER M1 ;
        RECT 9.904 23.652 9.936 24.396 ;
  LAYER M1 ;
        RECT 9.904 24.828 9.936 25.572 ;
  LAYER M1 ;
        RECT 9.904 26.004 9.936 26.748 ;
  LAYER M1 ;
        RECT 9.904 27.18 9.936 27.924 ;
  LAYER M1 ;
        RECT 9.904 28.356 9.936 29.1 ;
  LAYER M1 ;
        RECT 9.904 29.532 9.936 30.276 ;
  LAYER M1 ;
        RECT 10.064 22.476 10.096 23.22 ;
  LAYER M1 ;
        RECT 10.064 23.652 10.096 24.396 ;
  LAYER M1 ;
        RECT 10.064 24.828 10.096 25.572 ;
  LAYER M1 ;
        RECT 10.064 26.004 10.096 26.748 ;
  LAYER M1 ;
        RECT 10.064 27.18 10.096 27.924 ;
  LAYER M1 ;
        RECT 10.064 28.356 10.096 29.1 ;
  LAYER M1 ;
        RECT 10.064 29.532 10.096 30.276 ;
  LAYER M1 ;
        RECT 10.624 22.476 10.656 23.22 ;
  LAYER M1 ;
        RECT 10.624 23.316 10.656 23.556 ;
  LAYER M1 ;
        RECT 10.624 23.652 10.656 24.396 ;
  LAYER M1 ;
        RECT 10.624 24.492 10.656 24.732 ;
  LAYER M1 ;
        RECT 10.624 24.828 10.656 25.572 ;
  LAYER M1 ;
        RECT 10.624 25.668 10.656 25.908 ;
  LAYER M1 ;
        RECT 10.624 26.004 10.656 26.748 ;
  LAYER M1 ;
        RECT 10.624 26.844 10.656 27.084 ;
  LAYER M1 ;
        RECT 10.624 27.18 10.656 27.924 ;
  LAYER M1 ;
        RECT 10.624 28.02 10.656 28.26 ;
  LAYER M1 ;
        RECT 10.624 28.356 10.656 29.1 ;
  LAYER M1 ;
        RECT 10.624 29.196 10.656 29.436 ;
  LAYER M1 ;
        RECT 10.624 29.532 10.656 30.276 ;
  LAYER M1 ;
        RECT 10.624 30.372 10.656 30.612 ;
  LAYER M1 ;
        RECT 10.624 30.876 10.656 31.116 ;
  LAYER M1 ;
        RECT 10.544 22.476 10.576 23.22 ;
  LAYER M1 ;
        RECT 10.544 23.652 10.576 24.396 ;
  LAYER M1 ;
        RECT 10.544 24.828 10.576 25.572 ;
  LAYER M1 ;
        RECT 10.544 26.004 10.576 26.748 ;
  LAYER M1 ;
        RECT 10.544 27.18 10.576 27.924 ;
  LAYER M1 ;
        RECT 10.544 28.356 10.576 29.1 ;
  LAYER M1 ;
        RECT 10.544 29.532 10.576 30.276 ;
  LAYER M1 ;
        RECT 10.704 22.476 10.736 23.22 ;
  LAYER M1 ;
        RECT 10.704 23.652 10.736 24.396 ;
  LAYER M1 ;
        RECT 10.704 24.828 10.736 25.572 ;
  LAYER M1 ;
        RECT 10.704 26.004 10.736 26.748 ;
  LAYER M1 ;
        RECT 10.704 27.18 10.736 27.924 ;
  LAYER M1 ;
        RECT 10.704 28.356 10.736 29.1 ;
  LAYER M1 ;
        RECT 10.704 29.532 10.736 30.276 ;
  LAYER M1 ;
        RECT 11.264 22.476 11.296 23.22 ;
  LAYER M1 ;
        RECT 11.264 23.316 11.296 23.556 ;
  LAYER M1 ;
        RECT 11.264 23.652 11.296 24.396 ;
  LAYER M1 ;
        RECT 11.264 24.492 11.296 24.732 ;
  LAYER M1 ;
        RECT 11.264 24.828 11.296 25.572 ;
  LAYER M1 ;
        RECT 11.264 25.668 11.296 25.908 ;
  LAYER M1 ;
        RECT 11.264 26.004 11.296 26.748 ;
  LAYER M1 ;
        RECT 11.264 26.844 11.296 27.084 ;
  LAYER M1 ;
        RECT 11.264 27.18 11.296 27.924 ;
  LAYER M1 ;
        RECT 11.264 28.02 11.296 28.26 ;
  LAYER M1 ;
        RECT 11.264 28.356 11.296 29.1 ;
  LAYER M1 ;
        RECT 11.264 29.196 11.296 29.436 ;
  LAYER M1 ;
        RECT 11.264 29.532 11.296 30.276 ;
  LAYER M1 ;
        RECT 11.264 30.372 11.296 30.612 ;
  LAYER M1 ;
        RECT 11.264 30.876 11.296 31.116 ;
  LAYER M1 ;
        RECT 11.184 22.476 11.216 23.22 ;
  LAYER M1 ;
        RECT 11.184 23.652 11.216 24.396 ;
  LAYER M1 ;
        RECT 11.184 24.828 11.216 25.572 ;
  LAYER M1 ;
        RECT 11.184 26.004 11.216 26.748 ;
  LAYER M1 ;
        RECT 11.184 27.18 11.216 27.924 ;
  LAYER M1 ;
        RECT 11.184 28.356 11.216 29.1 ;
  LAYER M1 ;
        RECT 11.184 29.532 11.216 30.276 ;
  LAYER M1 ;
        RECT 11.344 22.476 11.376 23.22 ;
  LAYER M1 ;
        RECT 11.344 23.652 11.376 24.396 ;
  LAYER M1 ;
        RECT 11.344 24.828 11.376 25.572 ;
  LAYER M1 ;
        RECT 11.344 26.004 11.376 26.748 ;
  LAYER M1 ;
        RECT 11.344 27.18 11.376 27.924 ;
  LAYER M1 ;
        RECT 11.344 28.356 11.376 29.1 ;
  LAYER M1 ;
        RECT 11.344 29.532 11.376 30.276 ;
  LAYER M1 ;
        RECT 11.904 22.476 11.936 23.22 ;
  LAYER M1 ;
        RECT 11.904 23.316 11.936 23.556 ;
  LAYER M1 ;
        RECT 11.904 23.652 11.936 24.396 ;
  LAYER M1 ;
        RECT 11.904 24.492 11.936 24.732 ;
  LAYER M1 ;
        RECT 11.904 24.828 11.936 25.572 ;
  LAYER M1 ;
        RECT 11.904 25.668 11.936 25.908 ;
  LAYER M1 ;
        RECT 11.904 26.004 11.936 26.748 ;
  LAYER M1 ;
        RECT 11.904 26.844 11.936 27.084 ;
  LAYER M1 ;
        RECT 11.904 27.18 11.936 27.924 ;
  LAYER M1 ;
        RECT 11.904 28.02 11.936 28.26 ;
  LAYER M1 ;
        RECT 11.904 28.356 11.936 29.1 ;
  LAYER M1 ;
        RECT 11.904 29.196 11.936 29.436 ;
  LAYER M1 ;
        RECT 11.904 29.532 11.936 30.276 ;
  LAYER M1 ;
        RECT 11.904 30.372 11.936 30.612 ;
  LAYER M1 ;
        RECT 11.904 30.876 11.936 31.116 ;
  LAYER M1 ;
        RECT 11.824 22.476 11.856 23.22 ;
  LAYER M1 ;
        RECT 11.824 23.652 11.856 24.396 ;
  LAYER M1 ;
        RECT 11.824 24.828 11.856 25.572 ;
  LAYER M1 ;
        RECT 11.824 26.004 11.856 26.748 ;
  LAYER M1 ;
        RECT 11.824 27.18 11.856 27.924 ;
  LAYER M1 ;
        RECT 11.824 28.356 11.856 29.1 ;
  LAYER M1 ;
        RECT 11.824 29.532 11.856 30.276 ;
  LAYER M1 ;
        RECT 11.984 22.476 12.016 23.22 ;
  LAYER M1 ;
        RECT 11.984 23.652 12.016 24.396 ;
  LAYER M1 ;
        RECT 11.984 24.828 12.016 25.572 ;
  LAYER M1 ;
        RECT 11.984 26.004 12.016 26.748 ;
  LAYER M1 ;
        RECT 11.984 27.18 12.016 27.924 ;
  LAYER M1 ;
        RECT 11.984 28.356 12.016 29.1 ;
  LAYER M1 ;
        RECT 11.984 29.532 12.016 30.276 ;
  LAYER M1 ;
        RECT 12.544 22.476 12.576 23.22 ;
  LAYER M1 ;
        RECT 12.544 23.316 12.576 23.556 ;
  LAYER M1 ;
        RECT 12.544 23.652 12.576 24.396 ;
  LAYER M1 ;
        RECT 12.544 24.492 12.576 24.732 ;
  LAYER M1 ;
        RECT 12.544 24.828 12.576 25.572 ;
  LAYER M1 ;
        RECT 12.544 25.668 12.576 25.908 ;
  LAYER M1 ;
        RECT 12.544 26.004 12.576 26.748 ;
  LAYER M1 ;
        RECT 12.544 26.844 12.576 27.084 ;
  LAYER M1 ;
        RECT 12.544 27.18 12.576 27.924 ;
  LAYER M1 ;
        RECT 12.544 28.02 12.576 28.26 ;
  LAYER M1 ;
        RECT 12.544 28.356 12.576 29.1 ;
  LAYER M1 ;
        RECT 12.544 29.196 12.576 29.436 ;
  LAYER M1 ;
        RECT 12.544 29.532 12.576 30.276 ;
  LAYER M1 ;
        RECT 12.544 30.372 12.576 30.612 ;
  LAYER M1 ;
        RECT 12.544 30.876 12.576 31.116 ;
  LAYER M1 ;
        RECT 12.464 22.476 12.496 23.22 ;
  LAYER M1 ;
        RECT 12.464 23.652 12.496 24.396 ;
  LAYER M1 ;
        RECT 12.464 24.828 12.496 25.572 ;
  LAYER M1 ;
        RECT 12.464 26.004 12.496 26.748 ;
  LAYER M1 ;
        RECT 12.464 27.18 12.496 27.924 ;
  LAYER M1 ;
        RECT 12.464 28.356 12.496 29.1 ;
  LAYER M1 ;
        RECT 12.464 29.532 12.496 30.276 ;
  LAYER M1 ;
        RECT 12.624 22.476 12.656 23.22 ;
  LAYER M1 ;
        RECT 12.624 23.652 12.656 24.396 ;
  LAYER M1 ;
        RECT 12.624 24.828 12.656 25.572 ;
  LAYER M1 ;
        RECT 12.624 26.004 12.656 26.748 ;
  LAYER M1 ;
        RECT 12.624 27.18 12.656 27.924 ;
  LAYER M1 ;
        RECT 12.624 28.356 12.656 29.1 ;
  LAYER M1 ;
        RECT 12.624 29.532 12.656 30.276 ;
  LAYER M1 ;
        RECT 13.184 22.476 13.216 23.22 ;
  LAYER M1 ;
        RECT 13.184 23.316 13.216 23.556 ;
  LAYER M1 ;
        RECT 13.184 23.652 13.216 24.396 ;
  LAYER M1 ;
        RECT 13.184 24.492 13.216 24.732 ;
  LAYER M1 ;
        RECT 13.184 24.828 13.216 25.572 ;
  LAYER M1 ;
        RECT 13.184 25.668 13.216 25.908 ;
  LAYER M1 ;
        RECT 13.184 26.004 13.216 26.748 ;
  LAYER M1 ;
        RECT 13.184 26.844 13.216 27.084 ;
  LAYER M1 ;
        RECT 13.184 27.18 13.216 27.924 ;
  LAYER M1 ;
        RECT 13.184 28.02 13.216 28.26 ;
  LAYER M1 ;
        RECT 13.184 28.356 13.216 29.1 ;
  LAYER M1 ;
        RECT 13.184 29.196 13.216 29.436 ;
  LAYER M1 ;
        RECT 13.184 29.532 13.216 30.276 ;
  LAYER M1 ;
        RECT 13.184 30.372 13.216 30.612 ;
  LAYER M1 ;
        RECT 13.184 30.876 13.216 31.116 ;
  LAYER M1 ;
        RECT 13.104 22.476 13.136 23.22 ;
  LAYER M1 ;
        RECT 13.104 23.652 13.136 24.396 ;
  LAYER M1 ;
        RECT 13.104 24.828 13.136 25.572 ;
  LAYER M1 ;
        RECT 13.104 26.004 13.136 26.748 ;
  LAYER M1 ;
        RECT 13.104 27.18 13.136 27.924 ;
  LAYER M1 ;
        RECT 13.104 28.356 13.136 29.1 ;
  LAYER M1 ;
        RECT 13.104 29.532 13.136 30.276 ;
  LAYER M1 ;
        RECT 13.264 22.476 13.296 23.22 ;
  LAYER M1 ;
        RECT 13.264 23.652 13.296 24.396 ;
  LAYER M1 ;
        RECT 13.264 24.828 13.296 25.572 ;
  LAYER M1 ;
        RECT 13.264 26.004 13.296 26.748 ;
  LAYER M1 ;
        RECT 13.264 27.18 13.296 27.924 ;
  LAYER M1 ;
        RECT 13.264 28.356 13.296 29.1 ;
  LAYER M1 ;
        RECT 13.264 29.532 13.296 30.276 ;
  LAYER M1 ;
        RECT 13.824 22.476 13.856 23.22 ;
  LAYER M1 ;
        RECT 13.824 23.316 13.856 23.556 ;
  LAYER M1 ;
        RECT 13.824 23.652 13.856 24.396 ;
  LAYER M1 ;
        RECT 13.824 24.492 13.856 24.732 ;
  LAYER M1 ;
        RECT 13.824 24.828 13.856 25.572 ;
  LAYER M1 ;
        RECT 13.824 25.668 13.856 25.908 ;
  LAYER M1 ;
        RECT 13.824 26.004 13.856 26.748 ;
  LAYER M1 ;
        RECT 13.824 26.844 13.856 27.084 ;
  LAYER M1 ;
        RECT 13.824 27.18 13.856 27.924 ;
  LAYER M1 ;
        RECT 13.824 28.02 13.856 28.26 ;
  LAYER M1 ;
        RECT 13.824 28.356 13.856 29.1 ;
  LAYER M1 ;
        RECT 13.824 29.196 13.856 29.436 ;
  LAYER M1 ;
        RECT 13.824 29.532 13.856 30.276 ;
  LAYER M1 ;
        RECT 13.824 30.372 13.856 30.612 ;
  LAYER M1 ;
        RECT 13.824 30.876 13.856 31.116 ;
  LAYER M1 ;
        RECT 13.744 22.476 13.776 23.22 ;
  LAYER M1 ;
        RECT 13.744 23.652 13.776 24.396 ;
  LAYER M1 ;
        RECT 13.744 24.828 13.776 25.572 ;
  LAYER M1 ;
        RECT 13.744 26.004 13.776 26.748 ;
  LAYER M1 ;
        RECT 13.744 27.18 13.776 27.924 ;
  LAYER M1 ;
        RECT 13.744 28.356 13.776 29.1 ;
  LAYER M1 ;
        RECT 13.744 29.532 13.776 30.276 ;
  LAYER M1 ;
        RECT 13.904 22.476 13.936 23.22 ;
  LAYER M1 ;
        RECT 13.904 23.652 13.936 24.396 ;
  LAYER M1 ;
        RECT 13.904 24.828 13.936 25.572 ;
  LAYER M1 ;
        RECT 13.904 26.004 13.936 26.748 ;
  LAYER M1 ;
        RECT 13.904 27.18 13.936 27.924 ;
  LAYER M1 ;
        RECT 13.904 28.356 13.936 29.1 ;
  LAYER M1 ;
        RECT 13.904 29.532 13.936 30.276 ;
  LAYER M1 ;
        RECT 14.464 22.476 14.496 23.22 ;
  LAYER M1 ;
        RECT 14.464 23.316 14.496 23.556 ;
  LAYER M1 ;
        RECT 14.464 23.652 14.496 24.396 ;
  LAYER M1 ;
        RECT 14.464 24.492 14.496 24.732 ;
  LAYER M1 ;
        RECT 14.464 24.828 14.496 25.572 ;
  LAYER M1 ;
        RECT 14.464 25.668 14.496 25.908 ;
  LAYER M1 ;
        RECT 14.464 26.004 14.496 26.748 ;
  LAYER M1 ;
        RECT 14.464 26.844 14.496 27.084 ;
  LAYER M1 ;
        RECT 14.464 27.18 14.496 27.924 ;
  LAYER M1 ;
        RECT 14.464 28.02 14.496 28.26 ;
  LAYER M1 ;
        RECT 14.464 28.356 14.496 29.1 ;
  LAYER M1 ;
        RECT 14.464 29.196 14.496 29.436 ;
  LAYER M1 ;
        RECT 14.464 29.532 14.496 30.276 ;
  LAYER M1 ;
        RECT 14.464 30.372 14.496 30.612 ;
  LAYER M1 ;
        RECT 14.464 30.876 14.496 31.116 ;
  LAYER M1 ;
        RECT 14.384 22.476 14.416 23.22 ;
  LAYER M1 ;
        RECT 14.384 23.652 14.416 24.396 ;
  LAYER M1 ;
        RECT 14.384 24.828 14.416 25.572 ;
  LAYER M1 ;
        RECT 14.384 26.004 14.416 26.748 ;
  LAYER M1 ;
        RECT 14.384 27.18 14.416 27.924 ;
  LAYER M1 ;
        RECT 14.384 28.356 14.416 29.1 ;
  LAYER M1 ;
        RECT 14.384 29.532 14.416 30.276 ;
  LAYER M1 ;
        RECT 14.544 22.476 14.576 23.22 ;
  LAYER M1 ;
        RECT 14.544 23.652 14.576 24.396 ;
  LAYER M1 ;
        RECT 14.544 24.828 14.576 25.572 ;
  LAYER M1 ;
        RECT 14.544 26.004 14.576 26.748 ;
  LAYER M1 ;
        RECT 14.544 27.18 14.576 27.924 ;
  LAYER M1 ;
        RECT 14.544 28.356 14.576 29.1 ;
  LAYER M1 ;
        RECT 14.544 29.532 14.576 30.276 ;
  LAYER M1 ;
        RECT 15.104 22.476 15.136 23.22 ;
  LAYER M1 ;
        RECT 15.104 23.316 15.136 23.556 ;
  LAYER M1 ;
        RECT 15.104 23.652 15.136 24.396 ;
  LAYER M1 ;
        RECT 15.104 24.492 15.136 24.732 ;
  LAYER M1 ;
        RECT 15.104 24.828 15.136 25.572 ;
  LAYER M1 ;
        RECT 15.104 25.668 15.136 25.908 ;
  LAYER M1 ;
        RECT 15.104 26.004 15.136 26.748 ;
  LAYER M1 ;
        RECT 15.104 26.844 15.136 27.084 ;
  LAYER M1 ;
        RECT 15.104 27.18 15.136 27.924 ;
  LAYER M1 ;
        RECT 15.104 28.02 15.136 28.26 ;
  LAYER M1 ;
        RECT 15.104 28.356 15.136 29.1 ;
  LAYER M1 ;
        RECT 15.104 29.196 15.136 29.436 ;
  LAYER M1 ;
        RECT 15.104 29.532 15.136 30.276 ;
  LAYER M1 ;
        RECT 15.104 30.372 15.136 30.612 ;
  LAYER M1 ;
        RECT 15.104 30.876 15.136 31.116 ;
  LAYER M1 ;
        RECT 15.024 22.476 15.056 23.22 ;
  LAYER M1 ;
        RECT 15.024 23.652 15.056 24.396 ;
  LAYER M1 ;
        RECT 15.024 24.828 15.056 25.572 ;
  LAYER M1 ;
        RECT 15.024 26.004 15.056 26.748 ;
  LAYER M1 ;
        RECT 15.024 27.18 15.056 27.924 ;
  LAYER M1 ;
        RECT 15.024 28.356 15.056 29.1 ;
  LAYER M1 ;
        RECT 15.024 29.532 15.056 30.276 ;
  LAYER M1 ;
        RECT 15.184 22.476 15.216 23.22 ;
  LAYER M1 ;
        RECT 15.184 23.652 15.216 24.396 ;
  LAYER M1 ;
        RECT 15.184 24.828 15.216 25.572 ;
  LAYER M1 ;
        RECT 15.184 26.004 15.216 26.748 ;
  LAYER M1 ;
        RECT 15.184 27.18 15.216 27.924 ;
  LAYER M1 ;
        RECT 15.184 28.356 15.216 29.1 ;
  LAYER M1 ;
        RECT 15.184 29.532 15.216 30.276 ;
  LAYER M2 ;
        RECT 0.284 22.496 15.236 22.528 ;
  LAYER M2 ;
        RECT 0.924 22.58 14.596 22.612 ;
  LAYER M2 ;
        RECT 0.364 22.664 15.156 22.696 ;
  LAYER M2 ;
        RECT 0.364 23.336 15.156 23.368 ;
  LAYER M2 ;
        RECT 1.004 22.748 14.516 22.78 ;
  LAYER M2 ;
        RECT 0.924 23.672 14.596 23.704 ;
  LAYER M2 ;
        RECT 0.284 23.756 15.236 23.788 ;
  LAYER M2 ;
        RECT 1.004 23.84 14.516 23.872 ;
  LAYER M2 ;
        RECT 0.364 24.512 15.156 24.544 ;
  LAYER M2 ;
        RECT 0.364 23.924 15.156 23.956 ;
  LAYER M2 ;
        RECT 0.284 24.848 15.236 24.88 ;
  LAYER M2 ;
        RECT 0.924 24.932 14.596 24.964 ;
  LAYER M2 ;
        RECT 0.364 25.016 15.156 25.048 ;
  LAYER M2 ;
        RECT 0.364 25.688 15.156 25.72 ;
  LAYER M2 ;
        RECT 1.004 25.1 14.516 25.132 ;
  LAYER M2 ;
        RECT 0.924 26.024 14.596 26.056 ;
  LAYER M2 ;
        RECT 0.284 26.108 15.236 26.14 ;
  LAYER M2 ;
        RECT 1.004 26.192 14.516 26.224 ;
  LAYER M2 ;
        RECT 0.364 26.864 15.156 26.896 ;
  LAYER M2 ;
        RECT 0.364 26.276 15.156 26.308 ;
  LAYER M2 ;
        RECT 0.284 27.2 15.236 27.232 ;
  LAYER M2 ;
        RECT 0.924 27.284 14.596 27.316 ;
  LAYER M2 ;
        RECT 0.364 27.368 15.156 27.4 ;
  LAYER M2 ;
        RECT 0.364 28.04 15.156 28.072 ;
  LAYER M2 ;
        RECT 1.004 27.452 14.516 27.484 ;
  LAYER M2 ;
        RECT 0.924 28.376 14.596 28.408 ;
  LAYER M2 ;
        RECT 0.284 28.46 15.236 28.492 ;
  LAYER M2 ;
        RECT 1.004 28.544 14.516 28.576 ;
  LAYER M2 ;
        RECT 0.364 29.216 15.156 29.248 ;
  LAYER M2 ;
        RECT 0.364 28.628 15.156 28.66 ;
  LAYER M2 ;
        RECT 0.284 29.552 15.236 29.584 ;
  LAYER M2 ;
        RECT 0.924 29.636 14.596 29.668 ;
  LAYER M2 ;
        RECT 0.364 29.72 15.156 29.752 ;
  LAYER M2 ;
        RECT 0.364 30.392 15.156 30.424 ;
  LAYER M2 ;
        RECT 1.004 29.804 14.516 29.836 ;
  END 
END bandgap
