magic
tech scmos
timestamp 1597320842
<< nwell >>
rect -167 289 -115 347
rect -105 287 -63 347
rect -53 287 -17 347
rect -7 287 35 347
rect 45 287 87 347
rect 97 287 139 347
rect -47 281 -39 287
rect -7 -36 35 -5
rect 45 -36 87 -5
rect 97 -36 139 -5
<< psubstratepcontact >>
rect -160 -647 -149 -627
rect -136 -647 -125 -627
rect -113 -647 -102 -627
rect -91 -647 -80 -627
rect -70 -647 -59 -627
rect -49 -647 -38 -627
rect -27 -647 -16 -627
rect -5 -647 6 -627
rect 17 -647 28 -627
rect 38 -647 49 -627
rect 59 -647 70 -627
rect 79 -647 90 -627
rect 99 -647 110 -627
rect 119 -647 130 -627
rect 138 -647 149 -627
rect 158 -647 169 -627
rect 178 -647 189 -627
rect 199 -647 210 -627
rect 219 -647 230 -627
rect 240 -647 251 -627
rect 261 -647 272 -627
rect 280 -647 291 -627
rect 300 -647 311 -627
rect 320 -647 331 -627
rect 340 -647 351 -627
rect 359 -647 370 -627
rect 381 -647 392 -627
rect 404 -647 415 -627
rect 427 -647 438 -627
rect 450 -647 461 -627
rect 472 -647 483 -627
rect 494 -647 505 -627
rect 515 -647 526 -627
rect 535 -647 546 -627
<< nsubstratencontact >>
rect -164 321 -153 341
rect -146 321 -135 341
rect -129 321 -118 341
rect -102 321 -91 341
rect -77 321 -66 341
rect -50 321 -39 341
rect -31 321 -20 341
rect -4 321 7 341
rect 21 321 32 341
rect 48 321 59 341
rect 73 321 84 341
rect 100 321 111 341
rect 125 321 136 341
rect 149 321 160 341
rect 173 321 184 341
rect 195 321 206 341
rect 218 321 229 341
rect 240 321 251 341
rect 262 321 273 341
rect 285 321 296 341
rect 307 321 318 341
rect 329 321 340 341
rect 351 321 362 341
rect 374 321 385 341
rect 395 321 406 341
rect 416 321 427 341
rect 436 321 447 341
rect 457 321 468 341
rect 478 321 489 341
rect 499 321 510 341
rect 519 321 530 341
rect 536 321 547 341
rect 105 -385 125 -379
rect 105 -585 125 -579
rect 229 -391 249 -385
rect 445 -415 465 -409
<< polysilicon >>
rect -89 297 72 307
rect 80 297 123 307
rect -89 284 -79 297
rect 9 284 19 297
rect 61 284 71 297
rect 113 284 123 297
rect -146 191 -138 212
rect -39 150 -31 158
rect -70 142 -31 150
rect -72 -10 -69 -2
rect -33 -26 52 -16
rect 60 -26 123 -16
rect 9 -39 19 -26
rect 61 -39 71 -26
rect 113 -39 123 -26
rect -23 -353 0 -343
rect 8 -353 71 -343
rect -58 -366 -32 -358
rect 9 -366 19 -353
rect 61 -366 71 -353
<< polycontact >>
rect 72 297 80 307
rect -146 180 -138 191
rect -78 142 -70 150
rect -79 -10 -72 -2
rect -40 -26 -33 -16
rect 52 -26 60 -16
rect -30 -353 -23 -343
rect 0 -353 8 -343
rect -65 -366 -58 -358
<< metal1 >>
rect -167 321 -164 341
rect -153 321 -146 341
rect -135 321 -129 341
rect -118 321 -102 341
rect -91 321 -77 341
rect -66 321 -50 341
rect -39 321 -31 341
rect -20 321 -4 341
rect 7 321 21 341
rect 32 321 48 341
rect 59 321 73 341
rect 84 321 100 341
rect 111 321 125 341
rect 136 321 149 341
rect 160 321 173 341
rect 184 321 195 341
rect 206 321 218 341
rect 229 321 240 341
rect 251 321 262 341
rect 273 321 285 341
rect 296 321 307 341
rect 318 321 329 341
rect 340 321 351 341
rect 362 321 374 341
rect 385 321 395 341
rect 406 321 416 341
rect 427 321 436 341
rect 447 321 457 341
rect 468 321 478 341
rect 489 321 499 341
rect 510 321 519 341
rect 530 321 536 341
rect -160 281 -152 321
rect -98 281 -90 321
rect 0 284 8 321
rect 52 284 60 321
rect 72 284 80 297
rect 104 284 112 321
rect -160 -39 -152 215
rect -160 -627 -152 -49
rect -146 -65 -138 180
rect -130 -358 -122 215
rect -78 150 -70 161
rect -102 142 -78 150
rect -47 5 -40 161
rect -102 -39 -92 -17
rect -79 -65 -72 -10
rect -66 -26 -40 -16
rect -30 -343 -23 162
rect 20 -39 28 -2
rect 52 -39 60 -26
rect 72 -39 80 -2
rect 124 -39 132 -2
rect -130 -366 -65 -358
rect -30 -369 -23 -353
rect 0 -343 8 -325
rect 0 -366 8 -353
rect 52 -366 60 -325
rect 104 -345 112 -325
rect 104 -353 243 -345
rect 104 -379 197 -377
rect 104 -385 105 -379
rect 125 -385 197 -379
rect 235 -385 243 -353
rect -51 -627 -43 -445
rect 20 -599 28 -512
rect 72 -579 80 -512
rect 72 -585 105 -579
rect 327 -599 337 -339
rect 497 -409 507 -339
rect 465 -415 507 -409
rect 20 -607 337 -599
rect 538 -627 546 -312
rect -149 -647 -136 -627
rect -125 -647 -113 -627
rect -102 -647 -91 -627
rect -80 -647 -70 -627
rect -59 -647 -49 -627
rect -38 -647 -27 -627
rect -16 -647 -5 -627
rect 6 -647 17 -627
rect 28 -647 38 -627
rect 49 -647 59 -627
rect 70 -647 79 -627
rect 90 -647 99 -627
rect 110 -647 119 -627
rect 130 -647 138 -627
rect 149 -647 158 -627
rect 169 -647 178 -627
rect 189 -647 199 -627
rect 210 -647 219 -627
rect 230 -647 240 -627
rect 251 -647 261 -627
rect 272 -647 280 -627
rect 291 -647 300 -627
rect 311 -647 320 -627
rect 331 -647 340 -627
rect 351 -647 359 -627
rect 370 -647 381 -627
rect 392 -647 404 -627
rect 415 -647 427 -627
rect 438 -647 450 -627
rect 461 -647 472 -627
rect 483 -647 494 -627
rect 505 -647 515 -627
rect 526 -647 535 -627
<< m2contact >>
rect -160 -49 -152 -39
rect -146 -75 -138 -65
rect -102 -49 -92 -39
rect -79 -75 -72 -65
rect 327 -339 337 -329
rect 197 -385 207 -377
rect 497 -339 507 -329
<< metal2 >>
rect -152 -49 -102 -39
rect -138 -75 -79 -65
rect 197 -377 207 -322
rect 327 -329 337 -323
rect 497 -329 507 -313
<< pseudo_rnwell >>
rect 104 -379 126 -378
rect 104 -585 105 -379
rect 125 -585 126 -379
rect 104 -586 126 -585
rect 228 -385 250 -384
rect 228 -585 229 -385
rect 249 -564 250 -385
rect 255 -385 304 -384
rect 255 -564 256 -385
rect 249 -565 256 -564
rect 276 -406 283 -405
rect 276 -585 277 -406
rect 228 -586 277 -585
rect 282 -585 283 -406
rect 303 -564 304 -385
rect 309 -385 358 -384
rect 309 -564 310 -385
rect 303 -565 310 -564
rect 330 -406 337 -405
rect 330 -585 331 -406
rect 282 -586 331 -585
rect 336 -585 337 -406
rect 357 -564 358 -385
rect 363 -385 412 -384
rect 363 -564 364 -385
rect 357 -565 364 -564
rect 384 -406 391 -405
rect 384 -585 385 -406
rect 336 -586 385 -585
rect 390 -585 391 -406
rect 411 -564 412 -385
rect 417 -385 439 -384
rect 417 -564 418 -385
rect 411 -565 418 -564
rect 438 -564 439 -385
rect 444 -409 466 -408
rect 444 -564 445 -409
rect 438 -565 445 -564
rect 465 -585 466 -409
rect 390 -586 466 -585
<< rnwell >>
rect 105 -579 125 -385
rect 229 -565 249 -391
rect 256 -405 303 -385
rect 256 -565 276 -405
rect 229 -585 276 -565
rect 283 -565 303 -405
rect 310 -405 357 -385
rect 310 -565 330 -405
rect 283 -585 330 -565
rect 337 -565 357 -405
rect 364 -405 411 -385
rect 364 -565 384 -405
rect 337 -585 384 -565
rect 391 -565 411 -405
rect 418 -565 438 -385
rect 445 -565 465 -415
rect 391 -585 465 -565
use pd  pd_0
timestamp 1594499462
transform 1 0 -14 0 1 -429
box -38 -23 -8 63
use n1  n1_0
timestamp 1594253749
transform -1 0 28 0 1 -509
box -1 -3 29 143
use p1  p1_3
timestamp 1594254441
transform -1 0 19 0 1 -322
box -16 -6 26 286
use n1  n1_1
timestamp 1594253749
transform -1 0 80 0 1 -509
box -1 -3 29 143
use p1  p1_4
timestamp 1594254441
transform -1 0 71 0 1 -322
box -16 -6 26 286
use p1  p1_5
timestamp 1594254441
transform -1 0 123 0 1 -322
box -16 -6 26 286
use su3  su3_0
timestamp 1594543954
transform 1 0 -84 0 1 -98
box -28 72 -5 242
use pass  pass_0
timestamp 1594499169
transform 1 0 -65 0 -1 20
box -4 6 22 46
use p1  p1_0
timestamp 1594254441
transform 1 0 9 0 1 1
box -16 -6 26 286
use p1  p1_1
timestamp 1594254441
transform 1 0 61 0 1 1
box -16 -6 26 286
use p1  p1_2
timestamp 1594254441
transform 1 0 113 0 1 1
box -16 -6 26 286
use su1  su1_0
timestamp 1594254037
transform 1 0 -90 0 1 162
box -15 -7 27 125
use inv  inv_0
timestamp 1594513339
transform 1 0 -130 0 1 267
box -37 -55 15 22
use su2  su2_0
timestamp 1594254199
transform 1 0 -47 0 1 161
box -6 -6 30 126
use d1  d1_0
timestamp 1594590695
transform 0 -1 247 1 0 -313
box -10 -300 490 90
<< end >>
