magic
tech scmos
timestamp 1593520152
<< nwell >>
rect -11 0 1428 42
<< ntransistor >>
rect 361 -606 411 -586
rect 471 -606 521 -586
rect 581 -606 631 -586
rect 691 -606 741 -586
rect 801 -606 851 -586
rect 911 -606 961 -586
rect 1021 -606 1071 -586
rect 1131 -606 1181 -586
<< ptransistor >>
rect 55 6 105 36
rect 165 6 215 36
rect 275 6 325 36
rect 385 6 435 36
rect 495 6 545 36
rect 605 6 655 36
rect 715 6 765 36
rect 825 6 875 36
rect 935 6 985 36
rect 1045 6 1095 36
rect 1155 6 1205 36
rect 1265 6 1315 36
<< ndiffusion >>
rect 301 -606 361 -586
rect 411 -606 471 -586
rect 521 -606 581 -586
rect 631 -606 691 -586
rect 741 -606 801 -586
rect 851 -606 911 -586
rect 961 -606 1021 -586
rect 1071 -606 1131 -586
rect 1181 -606 1241 -586
<< pdiffusion >>
rect -5 26 55 36
rect -5 17 4 26
rect 11 17 16 26
rect 23 17 28 26
rect 35 17 40 26
rect 47 17 55 26
rect -5 6 55 17
rect 105 6 165 36
rect 215 26 275 36
rect 215 17 224 26
rect 231 17 236 26
rect 243 17 248 26
rect 255 17 259 26
rect 266 17 275 26
rect 215 6 275 17
rect 325 6 385 36
rect 435 26 495 36
rect 435 17 444 26
rect 451 17 456 26
rect 463 17 468 26
rect 475 17 479 26
rect 486 17 495 26
rect 435 6 495 17
rect 545 6 605 36
rect 655 27 715 36
rect 655 18 664 27
rect 671 18 676 27
rect 683 18 688 27
rect 695 18 699 27
rect 706 18 715 27
rect 655 6 715 18
rect 765 6 825 36
rect 875 27 935 36
rect 875 18 884 27
rect 891 18 896 27
rect 903 18 908 27
rect 915 18 919 27
rect 926 18 935 27
rect 875 6 935 18
rect 985 6 1045 36
rect 1095 27 1155 36
rect 1095 18 1104 27
rect 1111 18 1116 27
rect 1123 18 1128 27
rect 1135 18 1139 27
rect 1146 18 1155 27
rect 1095 6 1155 18
rect 1205 6 1265 36
rect 1315 27 1375 36
rect 1315 18 1324 27
rect 1331 18 1336 27
rect 1343 18 1348 27
rect 1355 18 1359 27
rect 1366 18 1375 27
rect 1315 6 1375 18
<< pdcontact >>
rect 4 17 11 26
rect 16 17 23 26
rect 28 17 35 26
rect 40 17 47 26
rect 224 17 231 26
rect 236 17 243 26
rect 248 17 255 26
rect 259 17 266 26
rect 444 17 451 26
rect 456 17 463 26
rect 468 17 475 26
rect 479 17 486 26
rect 664 18 671 27
rect 676 18 683 27
rect 688 18 695 27
rect 699 18 706 27
rect 884 18 891 27
rect 896 18 903 27
rect 908 18 915 27
rect 919 18 926 27
rect 1104 18 1111 27
rect 1116 18 1123 27
rect 1128 18 1135 27
rect 1139 18 1146 27
rect 1324 18 1331 27
rect 1336 18 1343 27
rect 1348 18 1355 27
rect 1359 18 1366 27
<< polysilicon >>
rect 72 69 1298 85
rect 72 39 88 69
rect 182 39 198 69
rect 292 39 308 69
rect 402 39 418 69
rect 512 39 528 69
rect 622 39 638 69
rect 732 39 748 69
rect 842 39 858 69
rect 952 39 968 69
rect 1062 39 1078 69
rect 1172 39 1188 69
rect 1282 39 1298 69
rect 55 36 105 39
rect 165 36 215 39
rect 275 36 325 39
rect 385 36 435 39
rect 495 36 545 39
rect 605 36 655 39
rect 715 36 765 39
rect 825 36 875 39
rect 935 36 985 39
rect 1045 36 1095 39
rect 1155 36 1205 39
rect 1265 36 1315 39
rect 55 3 105 6
rect 165 3 215 6
rect 275 3 325 6
rect 385 3 435 6
rect 495 3 545 6
rect 605 3 655 6
rect 715 3 765 6
rect 825 3 875 6
rect 935 3 985 6
rect 1045 3 1095 6
rect 1155 3 1205 6
rect 1265 3 1315 6
rect 378 -544 1164 -540
rect 378 -552 436 -544
rect 446 -552 876 -544
rect 886 -552 1164 -544
rect 378 -556 1164 -552
rect 378 -583 394 -556
rect 488 -583 504 -556
rect 598 -583 614 -556
rect 708 -583 724 -556
rect 818 -583 834 -556
rect 928 -583 944 -556
rect 1038 -583 1054 -556
rect 1148 -583 1164 -556
rect 361 -586 411 -583
rect 471 -586 521 -583
rect 581 -586 631 -583
rect 691 -586 741 -583
rect 801 -586 851 -583
rect 911 -586 961 -583
rect 1021 -586 1071 -583
rect 1131 -586 1181 -583
rect 361 -609 411 -606
rect 471 -609 521 -606
rect 581 -609 631 -606
rect 691 -609 741 -606
rect 801 -609 851 -606
rect 911 -609 961 -606
rect 1021 -609 1071 -606
rect 1131 -609 1181 -606
<< polycontact >>
rect 436 -552 446 -544
rect 876 -552 886 -544
<< metal1 >>
rect -17 101 1428 128
rect 15 32 35 101
rect 235 32 255 101
rect 455 32 475 101
rect 675 32 695 101
rect 895 32 915 101
rect 1115 32 1135 101
rect 1335 32 1355 101
rect 0 26 50 32
rect 0 17 4 26
rect 11 17 16 26
rect 23 17 28 26
rect 35 17 40 26
rect 47 17 50 26
rect 0 10 50 17
rect 110 10 160 32
rect 220 26 270 32
rect 220 17 224 26
rect 231 17 236 26
rect 243 17 248 26
rect 255 17 259 26
rect 266 17 270 26
rect 220 10 270 17
rect 330 10 380 32
rect 440 26 490 32
rect 440 17 444 26
rect 451 17 456 26
rect 463 17 468 26
rect 475 17 479 26
rect 486 17 490 26
rect 440 10 490 17
rect 550 10 600 32
rect 660 27 710 32
rect 660 18 664 27
rect 671 18 676 27
rect 683 18 688 27
rect 695 18 699 27
rect 706 18 710 27
rect 660 10 710 18
rect 770 10 820 32
rect 880 27 930 32
rect 880 18 884 27
rect 891 18 896 27
rect 903 18 908 27
rect 915 18 919 27
rect 926 18 930 27
rect 880 10 930 18
rect 990 10 1040 32
rect 1100 27 1150 32
rect 1100 18 1104 27
rect 1111 18 1116 27
rect 1123 18 1128 27
rect 1135 18 1139 27
rect 1146 18 1150 27
rect 1100 10 1150 18
rect 1210 10 1260 32
rect 1320 27 1370 32
rect 1320 18 1324 27
rect 1331 18 1336 27
rect 1343 18 1348 27
rect 1355 18 1359 27
rect 1366 18 1370 27
rect 1320 10 1370 18
rect 431 -524 891 -508
rect 431 -544 451 -524
rect 431 -552 436 -544
rect 446 -552 451 -544
rect 431 -588 451 -552
rect 871 -544 891 -524
rect 871 -552 876 -544
rect 886 -552 891 -544
rect 871 -588 891 -552
rect 306 -604 356 -588
rect 416 -604 466 -588
rect 526 -604 576 -588
rect 636 -604 686 -588
rect 746 -604 796 -588
rect 856 -604 906 -588
rect 966 -604 1016 -588
rect 1076 -604 1126 -588
rect 1186 -604 1236 -588
rect 651 -644 671 -604
rect 1091 -644 1111 -604
rect 651 -660 1111 -644
<< end >>
