* SPICE3 file created from new2.ext - technology: scmos

.option scale=0.1u

M1000 a_n213_118# a_n223_115# a_n243_118# w_n263_98# pfet w=80 l=10
+  ad=1600 pd=200 as=1600 ps=200
M1001 a_27_78# a_n23_75# a_n63_78# w_n83_58# pfet w=120 l=50
+  ad=4800 pd=320 as=4800 ps=320
M1002 a_377_n91# a_n23_n164# a_287_n91# w_n1073741817_n1073741817# nfet w=80 l=50
+  ad=3200 pd=240 as=3200 ps=240
M1003 a_547_78# a_n23_75# a_457_78# w_437_58# pfet w=120 l=50
+  ad=4800 pd=320 as=4800 ps=320
M1004 a_287_78# a_n23_75# a_197_78# w_177_58# pfet w=120 l=50
+  ad=4800 pd=320 as=4800 ps=320
M1005 a_27_n91# a_n23_n164# a_n63_n91# w_n1073741817_n1073741817# nfet w=80 l=50
+  ad=3200 pd=240 as=3200 ps=240
C0 a_n23_75# w_437_58# 2.01fF
C1 a_n23_75# w_177_58# 2.01fF
C2 a_n23_n164# w_n1073741817_n1073741817# 20.98fF
C3 a_n23_75# w_n1073741817_n1073741817# 30.50fF
C4 w_437_58# w_n1073741817_n1073741817# 20.67fF
C5 w_177_58# w_n1073741817_n1073741817# 20.67fF
C6 w_n83_58# w_n1073741817_n1073741817# 20.67fF
C7 w_n263_98# w_n1073741817_n1073741817# 8.21fF
C8 w_n523_78# w_n1073741817_n1073741817# 8.21fF **FLOATING
