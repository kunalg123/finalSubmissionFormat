* SPICE3 file created from su2.ext - technology: scmos

.option scale=0.1u

M1000 a_16_0# a_8_n3# a_0_0# w_n6_n6# pfet w=120 l=8
+  ad=960 pd=256 as=960 ps=256
C0 w_n6_n6# w_n1073741817_n1073741817# 3.61fF
