Bandgap reference with Start-Up

*Startup circuit
MSU1 3 2 1 1 p_mos W=3U L=0.2U
MSU2 3 3 4 4 n_mos W=0.2U L=0.2U
MSU3 4 4 5 5 n_mos W=0.2U L=0.2U
MSU4 5 5 0 0 n_mos W=0.2U L=0.2U
MSU5 8 3 7 7 p_mos W=3U L=0.2U
*................................
.ic   V(8)=0V V(9)=0V
M1 6 2 1 1 p_mos W=3U L=0.2U
M2 2 2 1 1 p_mos W=3U L=0.2U
M3 14 2 1 1 p_mos W=3U L=0.2U
M4 8 7 6 6 p_mos W=3U L=0.2U
M5 7 7 2 2 p_mos W=3U L=0.2U
M6 vref 7 14 14 p_mos W=3U L=0.2U
M7 8 8 9 9 n_mos W=1U L=0.2U
M8 7 8 11 11 n_mos W=1U L=0.2U
M9 9 9 10 10 n_mos W=1U L=0.2U
M10 11 9 12 12 n_mos W=1U L=0.2U
*................................
R1 12 13 2.2K
R2 vref 15 19K
D1 10 0 PNPDIODE
D2 13 0 PNPDIODE 8
D3 15 0 PNPDIODE 8
*................................
Vdd 1 0 dc 3.3
.model PNPDIODE D is=1e-18 n=1
.include osu018.lib
.tran 0.01 100ns
.control
run
plot v(vref) yl 0.6V 1.3V
.endc
.end
