* SPICE3 file created from m_l.ext - technology: scmos

.option scale=0.1u

M1000 a_n417_n20# a_n417_n20# b w_n1073741817_n1073741817# nfet w=30 l=10
+  ad=600 pd=100 as=600 ps=100
M1001 b b c w_n1073741817_n1073741817# nfet w=30 l=10
+  ad=0 pd=0 as=600 ps=100
M1002 c c a_n497_n17# w_n1073741817_n1073741817# nfet w=30 l=10
+  ad=0 pd=0 as=600 ps=100
