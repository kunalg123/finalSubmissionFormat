VBGP v/s Temperature [-40c - 140 ] 
M1 3 2 1 1 pfet W=wp L=ll
M2 2 2 1 1 pfet W=wp L=ll
M3 5 2 1 1 pfet W=wp L=ll


M4 6 4 3 1 pfet W=wp L=ll
M5 4 4 2 1 pfet W=wp L=ll
M6 vref 4 5 1 pfet W=wp L=ll


M7 6 6 7 0 nfet W=wn L=ll
M8 4 6 8 0 nfet W=wn L=ll



M9 a 2 1 1 pfet W=12U L=ll
M10 6 a 4 1 pfet W=12U L=0.8U
M11 a a b 0 nfet W=1U L=3u
M12 b b c 0 nfet W=1U L=3u
M13 c c 0 0 nfet W=1U L=3U


D1 7 0 PNPDIODE
R1 8 9 9K
D2 9 0 PNPDIODE 8
R2 vref 10 76K
D3 10 0 PNPDIODE 8
.param wp=28U wn=wp/2 ll=1U


Vdd 1 0 3.3
.model PNPDIODE D is=1e-18 n=1
.include osu018.lib
.dc temp -40 140 1
.control
run
plot v(vref)
.endc
.end
