magic
tech scmos
timestamp 1594286773
<< nsubstratencontact >>
rect 38 -487 58 -481
rect 280 -657 300 -650
<< pseudo_rnwell >>
rect 37 -481 59 -480
rect 37 -681 38 -481
rect 58 -660 59 -481
rect 67 -487 120 -486
rect 67 -660 68 -487
rect 58 -661 68 -660
rect 88 -508 99 -507
rect 88 -681 89 -508
rect 37 -682 89 -681
rect 98 -681 99 -508
rect 119 -660 120 -487
rect 128 -487 180 -486
rect 128 -660 129 -487
rect 119 -661 129 -660
rect 149 -508 159 -507
rect 149 -681 150 -508
rect 98 -682 150 -681
rect 158 -681 159 -508
rect 179 -660 180 -487
rect 188 -487 240 -486
rect 188 -660 189 -487
rect 179 -661 189 -660
rect 209 -508 219 -507
rect 209 -681 210 -508
rect 158 -682 210 -681
rect 218 -681 219 -508
rect 239 -660 240 -487
rect 248 -487 301 -486
rect 248 -660 249 -487
rect 239 -661 249 -660
rect 269 -508 280 -507
rect 269 -681 270 -508
rect 279 -657 280 -508
rect 300 -657 301 -487
rect 279 -658 301 -657
rect 218 -682 270 -681
<< rnwell >>
rect 38 -661 58 -487
rect 68 -507 119 -487
rect 68 -661 88 -507
rect 38 -681 88 -661
rect 99 -661 119 -507
rect 129 -507 179 -487
rect 129 -661 149 -507
rect 99 -681 149 -661
rect 159 -661 179 -507
rect 189 -507 239 -487
rect 189 -661 209 -507
rect 159 -681 209 -661
rect 219 -661 239 -507
rect 249 -507 300 -487
rect 249 -661 269 -507
rect 219 -681 269 -661
rect 280 -650 300 -507
<< labels >>
rlabel nsubstratencontact 290 -652 290 -652 1 b
rlabel nsubstratencontact 48 -484 48 -484 1 a
<< end >>
