* NGSPICE file created from bgr.ext - technology: scmos

.option scale=0.1u

M1000 3 2 1 1 pfet w=280 l=10
+  ad=5600 pd=1160 as=9600 ps=2000
M1001 2 2 1 1 pfet w=280 l=10
+  ad=5600 pd=1160 as=0 ps=0
M1002 5 2 1 1 pfet w=280 l=10
+  ad=5600 pd=1160 as=0 ps=0
M1003 6 4 3 1 pfet w=280 l=10
+  ad=3760 pd=836 as=0 ps=0
M1004 4 4 2 1 pfet w=280 l=10
+  ad=3760 pd=836 as=0 ps=0
M1005 vref 4 5 1 pfet w=280 l=10
+  ad=2800 pd=580 as=0 ps=0
M1006 6 6 7 0 nfet w=140 l=10
+  ad=1400 pd=300 as=1400 ps=300
M1007 4 6 8 0 nfet w=140 l=10
+  ad=1400 pd=300 as=1520 ps=352
M1008 a 2 1 1 pfet w=120 l=10
+  ad=1200 pd=260 as=0 ps=0
R0 vref 10 nwellResistor w=20 l=1637
M1009 a a m_l_0/b 0 nfet w=30 l=10
+  ad=600 pd=100 as=600 ps=100
M1010 m_l_0/b m_l_0/b m_l_0/c 0 nfet w=30 l=10
+  ad=0 pd=0 as=600 ps=100
M1011 m_l_0/c m_l_0/c 0 0 nfet w=30 l=10
+  ad=0 pd=0 as=600 ps=100
M1012 6 a 4 1 pfet w=120 l=8
+  ad=0 pd=0 as=0 ps=0
R1 9 8 nwellResistor w=20 l=194
C0 4 6 0.07fF
C1 10 r_0/a_37_n682# 0.02fF
C2 a 1 1.01fF
C3 vref r_0/a_37_n682# 0.02fF
C4 a m_l_0/b 0.04fF
C5 4 2 0.16fF
C6 m_l_0/b m_l_0/c 0.04fF
C7 1 3 0.43fF
C8 4 5 0.07fF
C9 6 1 0.36fF
C10 a 6 0.27fF
C11 vref 1 0.06fF
C12 4 1 3.42fF
C13 a 4 0.33fF
C14 2 1 5.59fF
C15 1 5 0.45fF
C16 4 3 0.07fF
C17 9 a_37_n688# 0.02fF
C18 8 a_37_n688# 0.02fF
C19 9 0 0.07fF
C20 a_37_n688# 0 2.95fF $ **FLOATING
C21 a 0 0.67fF
C22 m_l_0/b 0 0.55fF
C23 m_l_0/c 0 0.55fF
C24 vref 0 0.13fF
C25 r_0/a_37_n682# 0 27.31fF $ **FLOATING
C26 8 0 0.13fF
C27 7 0 0.20fF
C28 6 0 1.32fF
C29 4 0 1.59fF
C30 1 0 65.07fF
